MACRO INV_34777845_PG0
  ORIGIN 0 0 ;
  FOREIGN INV_34777845_PG0 0 0 ;
  SIZE 0.64 BY 4.704 ;
  PIN ZN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.124 2.252 0.356 2.284 ;
      LAYER M2 ;
        RECT 0.124 2.42 0.356 2.452 ;
      LAYER M2 ;
        RECT 0.124 2.252 0.196 2.284 ;
      LAYER M1 ;
        RECT 0.144 2.262 0.176 2.442 ;
      LAYER M2 ;
        RECT 0.124 2.42 0.196 2.452 ;
    END
  END ZN
  PIN I
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.124 1.412 0.356 1.444 ;
      LAYER M2 ;
        RECT 0.124 3.26 0.356 3.292 ;
      LAYER M2 ;
        RECT 0.124 1.412 0.196 1.444 ;
      LAYER M3 ;
        RECT 0.14 1.428 0.18 3.276 ;
      LAYER M2 ;
        RECT 0.124 3.26 0.196 3.292 ;
    END
  END I
  OBS 
  LAYER M1 ;
        RECT 0.304 1.56 0.336 2.304 ;
  LAYER M1 ;
        RECT 0.304 1.224 0.336 1.464 ;
  LAYER M1 ;
        RECT 0.304 0.468 0.336 0.708 ;
  LAYER M1 ;
        RECT 0.224 1.56 0.256 2.304 ;
  LAYER M1 ;
        RECT 0.384 1.56 0.416 2.304 ;
  LAYER M2 ;
        RECT 0.124 0.572 0.356 0.604 ;
  LAYER M2 ;
        RECT 0.204 2.168 0.436 2.2 ;
  LAYER M2 ;
        RECT 0.124 2.252 0.356 2.284 ;
  LAYER M2 ;
        RECT 0.124 1.412 0.356 1.444 ;
  LAYER M3 ;
        RECT 0.22 0.552 0.26 2.22 ;
  LAYER M1 ;
        RECT 0.304 2.4 0.336 3.144 ;
  LAYER M1 ;
        RECT 0.304 3.24 0.336 3.48 ;
  LAYER M1 ;
        RECT 0.304 3.996 0.336 4.236 ;
  LAYER M1 ;
        RECT 0.224 2.4 0.256 3.144 ;
  LAYER M1 ;
        RECT 0.384 2.4 0.416 3.144 ;
  LAYER M2 ;
        RECT 0.124 4.1 0.356 4.132 ;
  LAYER M2 ;
        RECT 0.204 2.504 0.436 2.536 ;
  LAYER M2 ;
        RECT 0.124 2.42 0.356 2.452 ;
  LAYER M2 ;
        RECT 0.124 3.26 0.356 3.292 ;
  LAYER M3 ;
        RECT 0.22 2.484 0.26 4.152 ;
  END 
END INV_34777845_PG0
