MACRO CCP_S_PMOS_B_12696969_X2_Y2
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CCP_S_PMOS_B_12696969_X2_Y2 0 0 ;
  SIZE 2560 BY 3528 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 2924 2276 2956 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1100 48 1140 2136 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1180 132 1220 2220 ;
    END
  END DB
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1260 216 1300 1464 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1340 300 1380 1548 ;
    END
  END SB
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1224 336 1968 ;
    LAYER M1 ;
      RECT 304 2064 336 2304 ;
    LAYER M1 ;
      RECT 304 2820 336 3060 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 224 1224 256 1968 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 384 1224 416 1968 ;
    LAYER M1 ;
      RECT 944 48 976 792 ;
    LAYER M1 ;
      RECT 944 888 976 1128 ;
    LAYER M1 ;
      RECT 944 1224 976 1968 ;
    LAYER M1 ;
      RECT 944 2064 976 2304 ;
    LAYER M1 ;
      RECT 944 2820 976 3060 ;
    LAYER M1 ;
      RECT 864 48 896 792 ;
    LAYER M1 ;
      RECT 864 1224 896 1968 ;
    LAYER M1 ;
      RECT 1024 48 1056 792 ;
    LAYER M1 ;
      RECT 1024 1224 1056 1968 ;
    LAYER M1 ;
      RECT 1584 48 1616 792 ;
    LAYER M1 ;
      RECT 1584 888 1616 1128 ;
    LAYER M1 ;
      RECT 1584 1224 1616 1968 ;
    LAYER M1 ;
      RECT 1584 2064 1616 2304 ;
    LAYER M1 ;
      RECT 1584 2820 1616 3060 ;
    LAYER M1 ;
      RECT 1504 48 1536 792 ;
    LAYER M1 ;
      RECT 1504 1224 1536 1968 ;
    LAYER M1 ;
      RECT 1664 48 1696 792 ;
    LAYER M1 ;
      RECT 1664 1224 1696 1968 ;
    LAYER M1 ;
      RECT 2224 48 2256 792 ;
    LAYER M1 ;
      RECT 2224 888 2256 1128 ;
    LAYER M1 ;
      RECT 2224 1224 2256 1968 ;
    LAYER M1 ;
      RECT 2224 2064 2256 2304 ;
    LAYER M1 ;
      RECT 2224 2820 2256 3060 ;
    LAYER M1 ;
      RECT 2144 48 2176 792 ;
    LAYER M1 ;
      RECT 2144 1224 2176 1968 ;
    LAYER M1 ;
      RECT 2304 48 2336 792 ;
    LAYER M1 ;
      RECT 2304 1224 2336 1968 ;
    LAYER M2 ;
      RECT 924 908 1636 940 ;
    LAYER M2 ;
      RECT 284 68 2276 100 ;
    LAYER M2 ;
      RECT 284 992 2276 1024 ;
    LAYER M2 ;
      RECT 924 152 1636 184 ;
    LAYER M2 ;
      RECT 204 236 2356 268 ;
    LAYER M2 ;
      RECT 844 320 1716 352 ;
    LAYER M2 ;
      RECT 284 2084 2276 2116 ;
    LAYER M2 ;
      RECT 924 1244 1636 1276 ;
    LAYER M2 ;
      RECT 924 2168 1636 2200 ;
    LAYER M2 ;
      RECT 284 1328 2276 1360 ;
    LAYER M2 ;
      RECT 844 1412 1716 1444 ;
    LAYER M2 ;
      RECT 204 1496 2356 1528 ;
    LAYER V1 ;
      RECT 1584 152 1616 184 ;
    LAYER V1 ;
      RECT 1584 908 1616 940 ;
    LAYER V1 ;
      RECT 1584 1244 1616 1276 ;
    LAYER V1 ;
      RECT 1584 2168 1616 2200 ;
    LAYER V1 ;
      RECT 1584 2924 1616 2956 ;
    LAYER V1 ;
      RECT 944 152 976 184 ;
    LAYER V1 ;
      RECT 944 908 976 940 ;
    LAYER V1 ;
      RECT 944 1244 976 1276 ;
    LAYER V1 ;
      RECT 944 2168 976 2200 ;
    LAYER V1 ;
      RECT 944 2924 976 2956 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 992 336 1024 ;
    LAYER V1 ;
      RECT 304 1328 336 1360 ;
    LAYER V1 ;
      RECT 304 2084 336 2116 ;
    LAYER V1 ;
      RECT 304 2924 336 2956 ;
    LAYER V1 ;
      RECT 2224 68 2256 100 ;
    LAYER V1 ;
      RECT 2224 992 2256 1024 ;
    LAYER V1 ;
      RECT 2224 1328 2256 1360 ;
    LAYER V1 ;
      RECT 2224 2084 2256 2116 ;
    LAYER V1 ;
      RECT 2224 2924 2256 2956 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 224 1496 256 1528 ;
    LAYER V1 ;
      RECT 2304 236 2336 268 ;
    LAYER V1 ;
      RECT 2304 1496 2336 1528 ;
    LAYER V1 ;
      RECT 2144 236 2176 268 ;
    LAYER V1 ;
      RECT 2144 1496 2176 1528 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 384 1496 416 1528 ;
    LAYER V1 ;
      RECT 864 320 896 352 ;
    LAYER V1 ;
      RECT 864 1412 896 1444 ;
    LAYER V1 ;
      RECT 1024 320 1056 352 ;
    LAYER V1 ;
      RECT 1024 1412 1056 1444 ;
    LAYER V1 ;
      RECT 1504 320 1536 352 ;
    LAYER V1 ;
      RECT 1504 1412 1536 1444 ;
    LAYER V1 ;
      RECT 1664 320 1696 352 ;
    LAYER V1 ;
      RECT 1664 1412 1696 1444 ;
    LAYER V2 ;
      RECT 1104 68 1136 100 ;
    LAYER V2 ;
      RECT 1104 908 1136 940 ;
    LAYER V2 ;
      RECT 1104 1244 1136 1276 ;
    LAYER V2 ;
      RECT 1104 2084 1136 2116 ;
    LAYER V2 ;
      RECT 1184 152 1216 184 ;
    LAYER V2 ;
      RECT 1184 992 1216 1024 ;
    LAYER V2 ;
      RECT 1184 1328 1216 1360 ;
    LAYER V2 ;
      RECT 1184 2168 1216 2200 ;
    LAYER V2 ;
      RECT 1264 236 1296 268 ;
    LAYER V2 ;
      RECT 1264 1412 1296 1444 ;
    LAYER V2 ;
      RECT 1344 320 1376 352 ;
    LAYER V2 ;
      RECT 1344 1496 1376 1528 ;
    LAYER V0 ;
      RECT 304 545 336 577 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1721 336 1753 ;
    LAYER V0 ;
      RECT 304 2084 336 2116 ;
    LAYER V0 ;
      RECT 304 2924 336 2956 ;
    LAYER V0 ;
      RECT 304 2924 336 2956 ;
    LAYER V0 ;
      RECT 224 545 256 577 ;
    LAYER V0 ;
      RECT 224 1721 256 1753 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 384 1721 416 1753 ;
    LAYER V0 ;
      RECT 944 545 976 577 ;
    LAYER V0 ;
      RECT 944 908 976 940 ;
    LAYER V0 ;
      RECT 944 1721 976 1753 ;
    LAYER V0 ;
      RECT 944 2084 976 2116 ;
    LAYER V0 ;
      RECT 944 2924 976 2956 ;
    LAYER V0 ;
      RECT 944 2924 976 2956 ;
    LAYER V0 ;
      RECT 864 545 896 577 ;
    LAYER V0 ;
      RECT 864 1721 896 1753 ;
    LAYER V0 ;
      RECT 1024 545 1056 577 ;
    LAYER V0 ;
      RECT 1024 1721 1056 1753 ;
    LAYER V0 ;
      RECT 1584 545 1616 577 ;
    LAYER V0 ;
      RECT 1584 908 1616 940 ;
    LAYER V0 ;
      RECT 1584 1721 1616 1753 ;
    LAYER V0 ;
      RECT 1584 2084 1616 2116 ;
    LAYER V0 ;
      RECT 1584 2924 1616 2956 ;
    LAYER V0 ;
      RECT 1584 2924 1616 2956 ;
    LAYER V0 ;
      RECT 1504 545 1536 577 ;
    LAYER V0 ;
      RECT 1504 1721 1536 1753 ;
    LAYER V0 ;
      RECT 1664 545 1696 577 ;
    LAYER V0 ;
      RECT 1664 1721 1696 1753 ;
    LAYER V0 ;
      RECT 2224 545 2256 577 ;
    LAYER V0 ;
      RECT 2224 908 2256 940 ;
    LAYER V0 ;
      RECT 2224 1721 2256 1753 ;
    LAYER V0 ;
      RECT 2224 2084 2256 2116 ;
    LAYER V0 ;
      RECT 2224 2924 2256 2956 ;
    LAYER V0 ;
      RECT 2224 2924 2256 2956 ;
    LAYER V0 ;
      RECT 2144 545 2176 577 ;
    LAYER V0 ;
      RECT 2144 1721 2176 1753 ;
    LAYER V0 ;
      RECT 2304 545 2336 577 ;
    LAYER V0 ;
      RECT 2304 1721 2336 1753 ;
  END
END CCP_S_PMOS_B_12696969_X2_Y2
