MACRO COMP_GM_STAGE_0415
  ORIGIN 0 0 ;
  FOREIGN COMP_GM_STAGE_0415 0 0 ;
  SIZE 2.612 BY 15.372 ;
  PIN OUTP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.524 4.604 0.756 4.636 ;
      LAYER M2 ;
        RECT 0.524 4.772 0.756 4.804 ;
      LAYER M2 ;
        RECT 0.524 4.604 0.596 4.636 ;
      LAYER M3 ;
        RECT 0.54 4.599 0.58 4.809 ;
      LAYER M2 ;
        RECT 0.524 4.772 0.596 4.804 ;
    END
  END OUTP
  PIN OUTM
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.804 4.604 2.036 4.636 ;
      LAYER M2 ;
        RECT 1.804 4.772 2.036 4.804 ;
      LAYER M2 ;
        RECT 1.804 4.604 1.876 4.636 ;
      LAYER M1 ;
        RECT 1.824 4.614 1.856 4.794 ;
      LAYER M2 ;
        RECT 1.804 4.772 1.876 4.804 ;
    END
  END OUTM
  PIN INP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.004 13.844 1.556 13.876 ;
    END
  END INP
  PIN INM
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.164 13.928 1.396 13.96 ;
    END
  END INM
  OBS 
  LAYER M3 ;
        RECT 1.02 1.392 1.06 2.304 ;
  LAYER M2 ;
        RECT 0.524 3.764 0.756 3.796 ;
  LAYER M2 ;
        RECT 0.524 5.612 0.756 5.644 ;
  LAYER M2 ;
        RECT 0.684 3.764 0.756 3.796 ;
  LAYER M1 ;
        RECT 0.704 3.78 0.736 5.628 ;
  LAYER M2 ;
        RECT 0.684 5.612 0.756 5.644 ;
  LAYER M2 ;
        RECT 1.004 6.956 1.236 6.988 ;
  LAYER M3 ;
        RECT 1.1 8.448 1.14 10.536 ;
  LAYER M3 ;
        RECT 1.02 2.268 1.06 3.78 ;
  LAYER M2 ;
        RECT 0.72 3.764 1.04 3.796 ;
  LAYER M2 ;
        RECT 0.684 5.612 0.756 5.644 ;
  LAYER M3 ;
        RECT 0.7 5.628 0.74 6.972 ;
  LAYER M2 ;
        RECT 0.72 6.956 1.04 6.988 ;
  LAYER M2 ;
        RECT 1.084 6.956 1.156 6.988 ;
  LAYER M3 ;
        RECT 1.1 6.972 1.14 8.484 ;
  LAYER M2 ;
        RECT 1.004 3.764 1.076 3.796 ;
  LAYER M3 ;
        RECT 1.02 3.744 1.06 3.816 ;
  LAYER M2 ;
        RECT 1.004 3.764 1.076 3.796 ;
  LAYER M3 ;
        RECT 1.02 3.744 1.06 3.816 ;
  LAYER M2 ;
        RECT 0.684 5.612 0.756 5.644 ;
  LAYER M3 ;
        RECT 0.7 5.592 0.74 5.664 ;
  LAYER M2 ;
        RECT 0.684 6.956 0.756 6.988 ;
  LAYER M3 ;
        RECT 0.7 6.936 0.74 7.008 ;
  LAYER M2 ;
        RECT 1.004 3.764 1.076 3.796 ;
  LAYER M3 ;
        RECT 1.02 3.744 1.06 3.816 ;
  LAYER M2 ;
        RECT 0.684 5.612 0.756 5.644 ;
  LAYER M3 ;
        RECT 0.7 5.592 0.74 5.664 ;
  LAYER M2 ;
        RECT 0.684 6.956 0.756 6.988 ;
  LAYER M3 ;
        RECT 0.7 6.936 0.74 7.008 ;
  LAYER M2 ;
        RECT 1.004 3.764 1.076 3.796 ;
  LAYER M3 ;
        RECT 1.02 3.744 1.06 3.816 ;
  LAYER M2 ;
        RECT 0.684 5.612 0.756 5.644 ;
  LAYER M3 ;
        RECT 0.7 5.592 0.74 5.664 ;
  LAYER M2 ;
        RECT 0.684 6.956 0.756 6.988 ;
  LAYER M3 ;
        RECT 0.7 6.936 0.74 7.008 ;
  LAYER M2 ;
        RECT 1.004 3.764 1.076 3.796 ;
  LAYER M3 ;
        RECT 1.02 3.744 1.06 3.816 ;
  LAYER M2 ;
        RECT 1.084 6.956 1.156 6.988 ;
  LAYER M3 ;
        RECT 1.1 6.936 1.14 7.008 ;
  LAYER M2 ;
        RECT 0.684 5.612 0.756 5.644 ;
  LAYER M3 ;
        RECT 0.7 5.592 0.74 5.664 ;
  LAYER M2 ;
        RECT 0.684 6.956 0.756 6.988 ;
  LAYER M3 ;
        RECT 0.7 6.936 0.74 7.008 ;
  LAYER M2 ;
        RECT 1.004 3.764 1.076 3.796 ;
  LAYER M3 ;
        RECT 1.02 3.744 1.06 3.816 ;
  LAYER M2 ;
        RECT 1.084 6.956 1.156 6.988 ;
  LAYER M3 ;
        RECT 1.1 6.936 1.14 7.008 ;
  LAYER M3 ;
        RECT 1.1 1.308 1.14 2.22 ;
  LAYER M2 ;
        RECT 1.804 3.764 2.036 3.796 ;
  LAYER M2 ;
        RECT 1.804 5.612 2.036 5.644 ;
  LAYER M2 ;
        RECT 1.804 3.764 1.876 3.796 ;
  LAYER M3 ;
        RECT 1.82 3.78 1.86 5.628 ;
  LAYER M2 ;
        RECT 1.804 5.612 1.876 5.644 ;
  LAYER M2 ;
        RECT 1.164 6.872 1.396 6.904 ;
  LAYER M3 ;
        RECT 1.18 8.364 1.22 10.452 ;
  LAYER M3 ;
        RECT 1.1 2.184 1.14 3.78 ;
  LAYER M4 ;
        RECT 1.12 3.76 1.84 3.8 ;
  LAYER M3 ;
        RECT 1.82 3.74 1.86 3.82 ;
  LAYER M2 ;
        RECT 1.804 5.612 1.876 5.644 ;
  LAYER M1 ;
        RECT 1.824 5.628 1.856 6.888 ;
  LAYER M2 ;
        RECT 1.36 6.872 1.84 6.904 ;
  LAYER M2 ;
        RECT 1.164 6.872 1.236 6.904 ;
  LAYER M3 ;
        RECT 1.18 6.888 1.22 8.4 ;
  LAYER M3 ;
        RECT 1.1 3.74 1.14 3.82 ;
  LAYER M4 ;
        RECT 1.08 3.76 1.16 3.8 ;
  LAYER M3 ;
        RECT 1.82 3.74 1.86 3.82 ;
  LAYER M4 ;
        RECT 1.8 3.76 1.88 3.8 ;
  LAYER M3 ;
        RECT 1.1 3.74 1.14 3.82 ;
  LAYER M4 ;
        RECT 1.08 3.76 1.16 3.8 ;
  LAYER M3 ;
        RECT 1.82 3.74 1.86 3.82 ;
  LAYER M4 ;
        RECT 1.8 3.76 1.88 3.8 ;
  LAYER M1 ;
        RECT 1.824 5.592 1.856 5.664 ;
  LAYER M2 ;
        RECT 1.804 5.612 1.876 5.644 ;
  LAYER M1 ;
        RECT 1.824 6.852 1.856 6.924 ;
  LAYER M2 ;
        RECT 1.804 6.872 1.876 6.904 ;
  LAYER M3 ;
        RECT 1.1 3.74 1.14 3.82 ;
  LAYER M4 ;
        RECT 1.08 3.76 1.16 3.8 ;
  LAYER M3 ;
        RECT 1.82 3.74 1.86 3.82 ;
  LAYER M4 ;
        RECT 1.8 3.76 1.88 3.8 ;
  LAYER M1 ;
        RECT 1.824 5.592 1.856 5.664 ;
  LAYER M2 ;
        RECT 1.804 5.612 1.876 5.644 ;
  LAYER M1 ;
        RECT 1.824 6.852 1.856 6.924 ;
  LAYER M2 ;
        RECT 1.804 6.872 1.876 6.904 ;
  LAYER M3 ;
        RECT 1.1 3.74 1.14 3.82 ;
  LAYER M4 ;
        RECT 1.08 3.76 1.16 3.8 ;
  LAYER M3 ;
        RECT 1.82 3.74 1.86 3.82 ;
  LAYER M4 ;
        RECT 1.8 3.76 1.88 3.8 ;
  LAYER M1 ;
        RECT 1.824 5.592 1.856 5.664 ;
  LAYER M2 ;
        RECT 1.804 5.612 1.876 5.644 ;
  LAYER M1 ;
        RECT 1.824 6.852 1.856 6.924 ;
  LAYER M2 ;
        RECT 1.804 6.872 1.876 6.904 ;
  LAYER M2 ;
        RECT 1.164 6.872 1.236 6.904 ;
  LAYER M3 ;
        RECT 1.18 6.852 1.22 6.924 ;
  LAYER M3 ;
        RECT 1.1 3.74 1.14 3.82 ;
  LAYER M4 ;
        RECT 1.08 3.76 1.16 3.8 ;
  LAYER M3 ;
        RECT 1.82 3.74 1.86 3.82 ;
  LAYER M4 ;
        RECT 1.8 3.76 1.88 3.8 ;
  LAYER M1 ;
        RECT 1.824 5.592 1.856 5.664 ;
  LAYER M2 ;
        RECT 1.804 5.612 1.876 5.644 ;
  LAYER M1 ;
        RECT 1.824 6.852 1.856 6.924 ;
  LAYER M2 ;
        RECT 1.804 6.872 1.876 6.904 ;
  LAYER M2 ;
        RECT 1.164 6.872 1.236 6.904 ;
  LAYER M3 ;
        RECT 1.18 6.852 1.22 6.924 ;
  LAYER M3 ;
        RECT 1.1 3.74 1.14 3.82 ;
  LAYER M4 ;
        RECT 1.08 3.76 1.16 3.8 ;
  LAYER M3 ;
        RECT 1.82 3.74 1.86 3.82 ;
  LAYER M4 ;
        RECT 1.8 3.76 1.88 3.8 ;
  LAYER M2 ;
        RECT 1.164 6.116 1.396 6.148 ;
  LAYER M2 ;
        RECT 1.164 11.492 1.396 11.524 ;
  LAYER M2 ;
        RECT 0.364 13.844 0.596 13.876 ;
  LAYER M2 ;
        RECT 1.36 6.116 1.44 6.148 ;
  LAYER M3 ;
        RECT 1.42 6.132 1.46 11.508 ;
  LAYER M2 ;
        RECT 1.36 11.492 1.44 11.524 ;
  LAYER M2 ;
        RECT 0.88 11.492 1.2 11.524 ;
  LAYER M1 ;
        RECT 0.864 11.508 0.896 13.86 ;
  LAYER M2 ;
        RECT 0.56 13.844 0.88 13.876 ;
  LAYER M2 ;
        RECT 1.404 6.116 1.476 6.148 ;
  LAYER M3 ;
        RECT 1.42 6.096 1.46 6.168 ;
  LAYER M2 ;
        RECT 1.404 11.492 1.476 11.524 ;
  LAYER M3 ;
        RECT 1.42 11.472 1.46 11.544 ;
  LAYER M2 ;
        RECT 1.404 6.116 1.476 6.148 ;
  LAYER M3 ;
        RECT 1.42 6.096 1.46 6.168 ;
  LAYER M2 ;
        RECT 1.404 11.492 1.476 11.524 ;
  LAYER M3 ;
        RECT 1.42 11.472 1.46 11.544 ;
  LAYER M1 ;
        RECT 0.864 11.472 0.896 11.544 ;
  LAYER M2 ;
        RECT 0.844 11.492 0.916 11.524 ;
  LAYER M1 ;
        RECT 0.864 13.824 0.896 13.896 ;
  LAYER M2 ;
        RECT 0.844 13.844 0.916 13.876 ;
  LAYER M2 ;
        RECT 1.404 6.116 1.476 6.148 ;
  LAYER M3 ;
        RECT 1.42 6.096 1.46 6.168 ;
  LAYER M2 ;
        RECT 1.404 11.492 1.476 11.524 ;
  LAYER M3 ;
        RECT 1.42 11.472 1.46 11.544 ;
  LAYER M1 ;
        RECT 0.864 11.472 0.896 11.544 ;
  LAYER M2 ;
        RECT 0.844 11.492 0.916 11.524 ;
  LAYER M1 ;
        RECT 0.864 13.824 0.896 13.896 ;
  LAYER M2 ;
        RECT 0.844 13.844 0.916 13.876 ;
  LAYER M2 ;
        RECT 1.404 6.116 1.476 6.148 ;
  LAYER M3 ;
        RECT 1.42 6.096 1.46 6.168 ;
  LAYER M2 ;
        RECT 1.404 11.492 1.476 11.524 ;
  LAYER M3 ;
        RECT 1.42 11.472 1.46 11.544 ;
  LAYER M2 ;
        RECT 1.004 10.652 1.236 10.684 ;
  LAYER M2 ;
        RECT 1.004 13.004 1.556 13.036 ;
  LAYER M3 ;
        RECT 1.26 9.12 1.3 10.368 ;
  LAYER M2 ;
        RECT 1.164 10.652 1.236 10.684 ;
  LAYER M3 ;
        RECT 1.18 10.668 1.22 13.02 ;
  LAYER M2 ;
        RECT 1.164 13.004 1.236 13.036 ;
  LAYER M2 ;
        RECT 1.2 10.652 1.28 10.684 ;
  LAYER M3 ;
        RECT 1.26 10.332 1.3 10.668 ;
  LAYER M2 ;
        RECT 1.164 10.652 1.236 10.684 ;
  LAYER M3 ;
        RECT 1.18 10.632 1.22 10.704 ;
  LAYER M2 ;
        RECT 1.164 13.004 1.236 13.036 ;
  LAYER M3 ;
        RECT 1.18 12.984 1.22 13.056 ;
  LAYER M2 ;
        RECT 1.164 10.652 1.236 10.684 ;
  LAYER M3 ;
        RECT 1.18 10.632 1.22 10.704 ;
  LAYER M2 ;
        RECT 1.164 13.004 1.236 13.036 ;
  LAYER M3 ;
        RECT 1.18 12.984 1.22 13.056 ;
  LAYER M2 ;
        RECT 1.164 10.652 1.236 10.684 ;
  LAYER M3 ;
        RECT 1.18 10.632 1.22 10.704 ;
  LAYER M2 ;
        RECT 1.164 13.004 1.236 13.036 ;
  LAYER M3 ;
        RECT 1.18 12.984 1.22 13.056 ;
  LAYER M2 ;
        RECT 1.244 10.652 1.316 10.684 ;
  LAYER M3 ;
        RECT 1.26 10.632 1.3 10.704 ;
  LAYER M2 ;
        RECT 1.164 10.652 1.236 10.684 ;
  LAYER M3 ;
        RECT 1.18 10.632 1.22 10.704 ;
  LAYER M2 ;
        RECT 1.164 13.004 1.236 13.036 ;
  LAYER M3 ;
        RECT 1.18 12.984 1.22 13.056 ;
  LAYER M2 ;
        RECT 1.244 10.652 1.316 10.684 ;
  LAYER M3 ;
        RECT 1.26 10.632 1.3 10.704 ;
  LAYER M2 ;
        RECT 1.164 10.736 1.396 10.768 ;
  LAYER M2 ;
        RECT 1.164 13.088 1.396 13.12 ;
  LAYER M3 ;
        RECT 1.34 9.036 1.38 10.284 ;
  LAYER M2 ;
        RECT 1.324 10.736 1.396 10.768 ;
  LAYER M3 ;
        RECT 1.34 10.752 1.38 13.104 ;
  LAYER M2 ;
        RECT 1.324 13.088 1.396 13.12 ;
  LAYER M3 ;
        RECT 1.34 10.248 1.38 10.752 ;
  LAYER M2 ;
        RECT 1.324 10.736 1.396 10.768 ;
  LAYER M3 ;
        RECT 1.34 10.716 1.38 10.788 ;
  LAYER M2 ;
        RECT 1.324 13.088 1.396 13.12 ;
  LAYER M3 ;
        RECT 1.34 13.068 1.38 13.14 ;
  LAYER M2 ;
        RECT 1.324 10.736 1.396 10.768 ;
  LAYER M3 ;
        RECT 1.34 10.716 1.38 10.788 ;
  LAYER M2 ;
        RECT 1.324 13.088 1.396 13.12 ;
  LAYER M3 ;
        RECT 1.34 13.068 1.38 13.14 ;
  LAYER M2 ;
        RECT 1.324 10.736 1.396 10.768 ;
  LAYER M3 ;
        RECT 1.34 10.716 1.38 10.788 ;
  LAYER M2 ;
        RECT 1.324 13.088 1.396 13.12 ;
  LAYER M3 ;
        RECT 1.34 13.068 1.38 13.14 ;
  LAYER M2 ;
        RECT 1.324 10.736 1.396 10.768 ;
  LAYER M3 ;
        RECT 1.34 10.716 1.38 10.788 ;
  LAYER M2 ;
        RECT 1.324 13.088 1.396 13.12 ;
  LAYER M3 ;
        RECT 1.34 13.068 1.38 13.14 ;
  LAYER M3 ;
        RECT 1.26 13.152 1.3 14.736 ;
  LAYER M2 ;
        RECT 0.364 13.004 0.596 13.036 ;
  LAYER M3 ;
        RECT 1.26 13.148 1.3 13.228 ;
  LAYER M4 ;
        RECT 0.88 13.168 1.28 13.208 ;
  LAYER M3 ;
        RECT 0.86 12.999 0.9 13.209 ;
  LAYER M2 ;
        RECT 0.56 13.004 0.88 13.036 ;
  LAYER M2 ;
        RECT 0.844 13.004 0.916 13.036 ;
  LAYER M3 ;
        RECT 0.86 12.984 0.9 13.056 ;
  LAYER M3 ;
        RECT 0.86 13.148 0.9 13.228 ;
  LAYER M4 ;
        RECT 0.84 13.168 0.92 13.208 ;
  LAYER M3 ;
        RECT 1.26 13.148 1.3 13.228 ;
  LAYER M4 ;
        RECT 1.24 13.168 1.32 13.208 ;
  LAYER M3 ;
        RECT 1.26 13.148 1.3 13.228 ;
  LAYER M4 ;
        RECT 1.24 13.168 1.32 13.208 ;
  LAYER M1 ;
        RECT 0.704 1.56 0.736 2.304 ;
  LAYER M1 ;
        RECT 0.704 1.224 0.736 1.464 ;
  LAYER M1 ;
        RECT 0.704 0.468 0.736 0.708 ;
  LAYER M1 ;
        RECT 0.624 1.56 0.656 2.304 ;
  LAYER M1 ;
        RECT 0.784 1.56 0.816 2.304 ;
  LAYER M1 ;
        RECT 0.864 1.56 0.896 2.304 ;
  LAYER M1 ;
        RECT 0.864 1.224 0.896 1.464 ;
  LAYER M1 ;
        RECT 0.864 0.468 0.896 0.708 ;
  LAYER M1 ;
        RECT 0.944 1.56 0.976 2.304 ;
  LAYER M1 ;
        RECT 1.024 1.56 1.056 2.304 ;
  LAYER M1 ;
        RECT 1.024 1.224 1.056 1.464 ;
  LAYER M1 ;
        RECT 1.024 0.468 1.056 0.708 ;
  LAYER M1 ;
        RECT 1.104 1.56 1.136 2.304 ;
  LAYER M1 ;
        RECT 1.184 1.56 1.216 2.304 ;
  LAYER M1 ;
        RECT 1.184 1.224 1.216 1.464 ;
  LAYER M1 ;
        RECT 1.184 0.468 1.216 0.708 ;
  LAYER M1 ;
        RECT 1.264 1.56 1.296 2.304 ;
  LAYER M1 ;
        RECT 1.344 1.56 1.376 2.304 ;
  LAYER M1 ;
        RECT 1.344 1.224 1.376 1.464 ;
  LAYER M1 ;
        RECT 1.344 0.468 1.376 0.708 ;
  LAYER M1 ;
        RECT 1.424 1.56 1.456 2.304 ;
  LAYER M1 ;
        RECT 1.504 1.56 1.536 2.304 ;
  LAYER M1 ;
        RECT 1.504 1.224 1.536 1.464 ;
  LAYER M1 ;
        RECT 1.504 0.468 1.536 0.708 ;
  LAYER M1 ;
        RECT 1.584 1.56 1.616 2.304 ;
  LAYER M1 ;
        RECT 1.664 1.56 1.696 2.304 ;
  LAYER M1 ;
        RECT 1.664 1.224 1.696 1.464 ;
  LAYER M1 ;
        RECT 1.664 0.468 1.696 0.708 ;
  LAYER M1 ;
        RECT 1.744 1.56 1.776 2.304 ;
  LAYER M1 ;
        RECT 1.824 1.56 1.856 2.304 ;
  LAYER M1 ;
        RECT 1.824 1.224 1.856 1.464 ;
  LAYER M1 ;
        RECT 1.824 0.468 1.856 0.708 ;
  LAYER M1 ;
        RECT 1.904 1.56 1.936 2.304 ;
  LAYER M2 ;
        RECT 0.844 1.412 1.716 1.444 ;
  LAYER M2 ;
        RECT 0.684 2.252 1.876 2.284 ;
  LAYER M2 ;
        RECT 0.684 1.328 1.876 1.36 ;
  LAYER M2 ;
        RECT 0.844 2.168 1.716 2.2 ;
  LAYER M2 ;
        RECT 0.684 0.572 1.876 0.604 ;
  LAYER M2 ;
        RECT 0.604 2.084 1.956 2.116 ;
  LAYER M3 ;
        RECT 1.02 1.392 1.06 2.304 ;
  LAYER M3 ;
        RECT 1.1 1.308 1.14 2.22 ;
  LAYER M3 ;
        RECT 1.18 0.552 1.22 2.136 ;
  LAYER M1 ;
        RECT 0.544 3.912 0.576 4.656 ;
  LAYER M1 ;
        RECT 0.544 3.576 0.576 3.816 ;
  LAYER M1 ;
        RECT 0.544 2.82 0.576 3.06 ;
  LAYER M1 ;
        RECT 0.624 3.912 0.656 4.656 ;
  LAYER M1 ;
        RECT 0.464 3.912 0.496 4.656 ;
  LAYER M2 ;
        RECT 0.524 2.924 0.756 2.956 ;
  LAYER M2 ;
        RECT 0.444 4.52 0.676 4.552 ;
  LAYER M2 ;
        RECT 0.524 4.604 0.756 4.636 ;
  LAYER M2 ;
        RECT 0.524 3.764 0.756 3.796 ;
  LAYER M3 ;
        RECT 0.62 2.904 0.66 4.572 ;
  LAYER M1 ;
        RECT 0.544 4.752 0.576 5.496 ;
  LAYER M1 ;
        RECT 0.544 5.592 0.576 5.832 ;
  LAYER M1 ;
        RECT 0.544 6.348 0.576 6.588 ;
  LAYER M1 ;
        RECT 0.624 4.752 0.656 5.496 ;
  LAYER M1 ;
        RECT 0.464 4.752 0.496 5.496 ;
  LAYER M2 ;
        RECT 0.524 6.452 0.756 6.484 ;
  LAYER M2 ;
        RECT 0.444 4.856 0.676 4.888 ;
  LAYER M2 ;
        RECT 0.524 4.772 0.756 4.804 ;
  LAYER M2 ;
        RECT 0.524 5.612 0.756 5.644 ;
  LAYER M3 ;
        RECT 0.62 4.836 0.66 6.504 ;
  LAYER M1 ;
        RECT 1.984 3.912 2.016 4.656 ;
  LAYER M1 ;
        RECT 1.984 3.576 2.016 3.816 ;
  LAYER M1 ;
        RECT 1.984 2.82 2.016 3.06 ;
  LAYER M1 ;
        RECT 1.904 3.912 1.936 4.656 ;
  LAYER M1 ;
        RECT 2.064 3.912 2.096 4.656 ;
  LAYER M2 ;
        RECT 1.804 2.924 2.036 2.956 ;
  LAYER M2 ;
        RECT 1.884 4.52 2.116 4.552 ;
  LAYER M2 ;
        RECT 1.804 4.604 2.036 4.636 ;
  LAYER M2 ;
        RECT 1.804 3.764 2.036 3.796 ;
  LAYER M3 ;
        RECT 1.9 2.904 1.94 4.572 ;
  LAYER M1 ;
        RECT 1.984 4.752 2.016 5.496 ;
  LAYER M1 ;
        RECT 1.984 5.592 2.016 5.832 ;
  LAYER M1 ;
        RECT 1.984 6.348 2.016 6.588 ;
  LAYER M1 ;
        RECT 1.904 4.752 1.936 5.496 ;
  LAYER M1 ;
        RECT 2.064 4.752 2.096 5.496 ;
  LAYER M2 ;
        RECT 1.804 6.452 2.036 6.484 ;
  LAYER M2 ;
        RECT 1.884 4.856 2.116 4.888 ;
  LAYER M2 ;
        RECT 1.804 4.772 2.036 4.804 ;
  LAYER M2 ;
        RECT 1.804 5.612 2.036 5.644 ;
  LAYER M3 ;
        RECT 1.9 4.836 1.94 6.504 ;
  LAYER M1 ;
        RECT 1.184 6.264 1.216 7.008 ;
  LAYER M1 ;
        RECT 1.184 5.928 1.216 6.168 ;
  LAYER M1 ;
        RECT 1.184 5.172 1.216 5.412 ;
  LAYER M1 ;
        RECT 1.104 6.264 1.136 7.008 ;
  LAYER M1 ;
        RECT 1.264 6.264 1.296 7.008 ;
  LAYER M1 ;
        RECT 1.344 6.264 1.376 7.008 ;
  LAYER M1 ;
        RECT 1.344 5.928 1.376 6.168 ;
  LAYER M1 ;
        RECT 1.344 5.172 1.376 5.412 ;
  LAYER M1 ;
        RECT 1.424 6.264 1.456 7.008 ;
  LAYER M2 ;
        RECT 1.164 5.276 1.396 5.308 ;
  LAYER M2 ;
        RECT 1.084 6.788 1.476 6.82 ;
  LAYER M2 ;
        RECT 1.004 6.956 1.236 6.988 ;
  LAYER M2 ;
        RECT 1.164 6.872 1.396 6.904 ;
  LAYER M2 ;
        RECT 1.164 6.116 1.396 6.148 ;
  LAYER M3 ;
        RECT 1.26 5.256 1.3 6.84 ;
  LAYER M1 ;
        RECT 1.184 10.632 1.216 11.376 ;
  LAYER M1 ;
        RECT 1.184 11.472 1.216 11.712 ;
  LAYER M1 ;
        RECT 1.184 12.228 1.216 12.468 ;
  LAYER M1 ;
        RECT 1.104 10.632 1.136 11.376 ;
  LAYER M1 ;
        RECT 1.264 10.632 1.296 11.376 ;
  LAYER M1 ;
        RECT 1.344 10.632 1.376 11.376 ;
  LAYER M1 ;
        RECT 1.344 11.472 1.376 11.712 ;
  LAYER M1 ;
        RECT 1.344 12.228 1.376 12.468 ;
  LAYER M1 ;
        RECT 1.424 10.632 1.456 11.376 ;
  LAYER M2 ;
        RECT 1.164 12.332 1.396 12.364 ;
  LAYER M2 ;
        RECT 1.084 10.82 1.476 10.852 ;
  LAYER M2 ;
        RECT 1.004 10.652 1.236 10.684 ;
  LAYER M2 ;
        RECT 1.164 10.736 1.396 10.768 ;
  LAYER M2 ;
        RECT 1.164 11.492 1.396 11.524 ;
  LAYER M3 ;
        RECT 1.26 10.8 1.3 12.384 ;
  LAYER M1 ;
        RECT 1.024 12.984 1.056 13.728 ;
  LAYER M1 ;
        RECT 1.024 13.824 1.056 14.064 ;
  LAYER M1 ;
        RECT 1.024 14.58 1.056 14.82 ;
  LAYER M1 ;
        RECT 0.944 12.984 0.976 13.728 ;
  LAYER M1 ;
        RECT 1.104 12.984 1.136 13.728 ;
  LAYER M1 ;
        RECT 1.184 12.984 1.216 13.728 ;
  LAYER M1 ;
        RECT 1.184 13.824 1.216 14.064 ;
  LAYER M1 ;
        RECT 1.184 14.58 1.216 14.82 ;
  LAYER M1 ;
        RECT 1.264 12.984 1.296 13.728 ;
  LAYER M1 ;
        RECT 1.344 12.984 1.376 13.728 ;
  LAYER M1 ;
        RECT 1.344 13.824 1.376 14.064 ;
  LAYER M1 ;
        RECT 1.344 14.58 1.376 14.82 ;
  LAYER M1 ;
        RECT 1.424 12.984 1.456 13.728 ;
  LAYER M1 ;
        RECT 1.504 12.984 1.536 13.728 ;
  LAYER M1 ;
        RECT 1.504 13.824 1.536 14.064 ;
  LAYER M1 ;
        RECT 1.504 14.58 1.536 14.82 ;
  LAYER M1 ;
        RECT 1.584 12.984 1.616 13.728 ;
  LAYER M2 ;
        RECT 1.004 14.684 1.556 14.716 ;
  LAYER M2 ;
        RECT 0.924 13.172 1.636 13.204 ;
  LAYER M2 ;
        RECT 1.004 13.004 1.556 13.036 ;
  LAYER M2 ;
        RECT 1.164 13.088 1.396 13.12 ;
  LAYER M2 ;
        RECT 1.004 13.844 1.556 13.876 ;
  LAYER M2 ;
        RECT 1.164 13.928 1.396 13.96 ;
  LAYER M3 ;
        RECT 1.26 13.152 1.3 14.736 ;
  LAYER M1 ;
        RECT 0.304 9.792 0.336 10.536 ;
  LAYER M1 ;
        RECT 0.304 9.456 0.336 9.696 ;
  LAYER M1 ;
        RECT 0.304 8.616 0.336 9.36 ;
  LAYER M1 ;
        RECT 0.304 8.28 0.336 8.52 ;
  LAYER M1 ;
        RECT 0.304 7.524 0.336 7.764 ;
  LAYER M1 ;
        RECT 0.224 9.792 0.256 10.536 ;
  LAYER M1 ;
        RECT 0.224 8.616 0.256 9.36 ;
  LAYER M1 ;
        RECT 0.384 9.792 0.416 10.536 ;
  LAYER M1 ;
        RECT 0.384 8.616 0.416 9.36 ;
  LAYER M1 ;
        RECT 0.944 9.792 0.976 10.536 ;
  LAYER M1 ;
        RECT 0.944 9.456 0.976 9.696 ;
  LAYER M1 ;
        RECT 0.944 8.616 0.976 9.36 ;
  LAYER M1 ;
        RECT 0.944 8.28 0.976 8.52 ;
  LAYER M1 ;
        RECT 0.944 7.524 0.976 7.764 ;
  LAYER M1 ;
        RECT 0.864 9.792 0.896 10.536 ;
  LAYER M1 ;
        RECT 0.864 8.616 0.896 9.36 ;
  LAYER M1 ;
        RECT 1.024 9.792 1.056 10.536 ;
  LAYER M1 ;
        RECT 1.024 8.616 1.056 9.36 ;
  LAYER M1 ;
        RECT 1.584 9.792 1.616 10.536 ;
  LAYER M1 ;
        RECT 1.584 9.456 1.616 9.696 ;
  LAYER M1 ;
        RECT 1.584 8.616 1.616 9.36 ;
  LAYER M1 ;
        RECT 1.584 8.28 1.616 8.52 ;
  LAYER M1 ;
        RECT 1.584 7.524 1.616 7.764 ;
  LAYER M1 ;
        RECT 1.504 9.792 1.536 10.536 ;
  LAYER M1 ;
        RECT 1.504 8.616 1.536 9.36 ;
  LAYER M1 ;
        RECT 1.664 9.792 1.696 10.536 ;
  LAYER M1 ;
        RECT 1.664 8.616 1.696 9.36 ;
  LAYER M1 ;
        RECT 2.224 9.792 2.256 10.536 ;
  LAYER M1 ;
        RECT 2.224 9.456 2.256 9.696 ;
  LAYER M1 ;
        RECT 2.224 8.616 2.256 9.36 ;
  LAYER M1 ;
        RECT 2.224 8.28 2.256 8.52 ;
  LAYER M1 ;
        RECT 2.224 7.524 2.256 7.764 ;
  LAYER M1 ;
        RECT 2.144 9.792 2.176 10.536 ;
  LAYER M1 ;
        RECT 2.144 8.616 2.176 9.36 ;
  LAYER M1 ;
        RECT 2.304 9.792 2.336 10.536 ;
  LAYER M1 ;
        RECT 2.304 8.616 2.336 9.36 ;
  LAYER M2 ;
        RECT 0.924 9.644 1.636 9.676 ;
  LAYER M2 ;
        RECT 0.284 10.484 2.276 10.516 ;
  LAYER M2 ;
        RECT 0.284 9.56 2.276 9.592 ;
  LAYER M2 ;
        RECT 0.924 10.4 1.636 10.432 ;
  LAYER M2 ;
        RECT 0.204 10.316 2.356 10.348 ;
  LAYER M2 ;
        RECT 0.844 10.232 1.716 10.264 ;
  LAYER M2 ;
        RECT 0.284 8.468 2.276 8.5 ;
  LAYER M2 ;
        RECT 0.924 9.308 1.636 9.34 ;
  LAYER M2 ;
        RECT 0.924 8.384 1.636 8.416 ;
  LAYER M2 ;
        RECT 0.284 9.224 2.276 9.256 ;
  LAYER M2 ;
        RECT 0.844 9.14 1.716 9.172 ;
  LAYER M2 ;
        RECT 0.204 9.056 2.356 9.088 ;
  LAYER M2 ;
        RECT 0.284 7.628 2.276 7.66 ;
  LAYER M3 ;
        RECT 1.1 8.448 1.14 10.536 ;
  LAYER M3 ;
        RECT 1.18 8.364 1.22 10.452 ;
  LAYER M3 ;
        RECT 1.26 9.12 1.3 10.368 ;
  LAYER M3 ;
        RECT 1.34 9.036 1.38 10.284 ;
  LAYER M1 ;
        RECT 0.384 12.984 0.416 13.728 ;
  LAYER M1 ;
        RECT 0.384 13.824 0.416 14.064 ;
  LAYER M1 ;
        RECT 0.384 14.58 0.416 14.82 ;
  LAYER M1 ;
        RECT 0.464 12.984 0.496 13.728 ;
  LAYER M1 ;
        RECT 0.304 12.984 0.336 13.728 ;
  LAYER M2 ;
        RECT 0.364 14.684 0.596 14.716 ;
  LAYER M2 ;
        RECT 0.284 13.088 0.516 13.12 ;
  LAYER M2 ;
        RECT 0.364 13.004 0.596 13.036 ;
  LAYER M2 ;
        RECT 0.364 13.844 0.596 13.876 ;
  LAYER M3 ;
        RECT 0.46 13.068 0.5 14.736 ;
  END 
END COMP_GM_STAGE_0415
