.subckt BUFFER_VREFP_ud GND IBIAS1 IBIAS2 VDD VREF VREFP VBK_1 VBK_2 VFB_IN VFB_O
M60  VREFP VREFP VREFP VDD pfet w=2u l=100n nf=4 nfin=4
M37  VDD net057 VDD VDD pfet w=5u l=5u nf=2 nfin=4
M29  VBK_2 net057 VREFP VDD pfet w=3u l=100n nf=6 nfin=4
M27  net057 net057 VFB_O VDD pfet w=0.25u l=100n nf=2 nfin=4
M28  VREFP VBK_1 VDD VDD pfet w=2.55u l=100n nf=6 nfin=4
M15  VFB_O net036 VDD VDD pfet w=212.5n l=100n nf=2 nfin=4
M59  net057 net057 net057 VDD pfet w=1u l=100n nf=2 nfin=4
M58  VFB_O VFB_O VFB_O VDD pfet w=1u l=100n nf=2 nfin=4
M54  VFB_O VFB_O VFB_O VDD pfet w=0.85u l=100n nf=2 nfin=4
M38  VDD net036 VDD VDD pfet w=0.5u l=2u nf=2 nfin=4
M65  IBIAS2 IBIAS2 IBIAS2 GND nfet w=150n l=100n nf=2 nfin=4
M64  IBIAS2 IBIAS2 GND GND nfet w=37.5n l=100n nf=2 nfin=4
M56  net057 net057 net057 GND nfet w=150n l=100n nf=2 nfin=4
M30  VBK_2 IBIAS2 GND GND nfet w=450n l=100n nf=6 nfin=4
M21  net057 IBIAS2 GND GND nfet w=37.5n l=100n nf=2 nfin=4
M12  net051 VREF net212 GND nfet w=50n l=100n nf=2 nfin=4
M11  net211 VREF net212 GND nfet w=50n l=100n nf=2 nfin=4
M10  net054 VFB_IN net212 GND nfet w=50n l=100n nf=2 nfin=4
M8  net215 VFB_IN net212 GND nfet w=50n l=100n nf=2 nfin=4
M5  net204 IBIAS1 GND GND nfet w=37.5n l=100n nf=2 nfin=4
M4  IBIAS1 IBIAS1 GND GND nfet w=37.5n l=100n nf=2 nfin=4
M3  net212 IBIAS1 GND GND nfet w=300n l=100n nf=4 nfin=4
M1  net207 net207 GND GND nfet w=37.5n l=650.0n nf=2 nfin=4
M6  net036 net207 GND GND nfet w=37.5n l=650.0n nf=2 nfin=4
M43  net211 net211 net211 GND nfet w=200n l=100n nf=2 nfin=4
M52  net036 net036 net036 GND nfet w=37.5n l=650.0n nf=2 nfin=4
M47  net212 net212 net212 GND nfet w=200n l=100n nf=2 nfin=4
M50  net207 net207 net207 GND nfet w=37.5n l=650.0n nf=2 nfin=4
M45  net051 net051 net051 GND nfet w=200n l=100n nf=2 nfin=4
M48  net212 net212 net212 GND nfet w=200n l=100n nf=2 nfin=4
M40  net204 net204 net204 GND nfet w=150n l=100n nf=2 nfin=4
M46  net054 net054 net054 GND nfet w=200n l=100n nf=2 nfin=4
M44  net215 net215 net215 GND nfet w=200n l=100n nf=2 nfin=4
M39  IBIAS1 IBIAS1 IBIAS1 GND nfet w=150n l=100n nf=2 nfin=4
M42  net051 net051 net051 VDD pfet w=0.6u l=100n nf=4 nfin=4
M35  net211 net211 net211 VDD pfet w=400n l=100n nf=2 nfin=4
M26  net054 net211 VDD VDD pfet w=0.8u l=100n nf=4 nfin=4
M25  net211 net211 VDD VDD pfet w=100n l=100n nf=2 nfin=4
M24  net051 net215 VDD VDD pfet w=0.8u l=100n nf=4 nfin=4
M23  net215 net215 VDD VDD pfet w=100n l=100n nf=2 nfin=4
M22  net204 net204 VDD VDD pfet w=125n l=500n nf=2 nfin=4
M41  net054 net054 net054 VDD pfet w=0.6u l=100n nf=4 nfin=4
M14  net207 net204 net054 VDD pfet w=300n l=100n nf=2 nfin=4
M13  net036 net204 net051 VDD pfet w=300n l=100n nf=2 nfin=4
M36  net215 net215 net215 VDD pfet w=400n l=100n nf=2 nfin=4
M31  net204 net204 net204 VDD pfet w=125n l=500n nf=2 nfin=4
.ends BUFFER_VREFP_ud

