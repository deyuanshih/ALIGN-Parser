MACRO SCM_NMOS_57551371
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_57551371 0 0 ;
  SIZE 1440 BY 2352 ;
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 460 48 500 960 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 152 1156 184 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 620 216 660 1800 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1644 336 1884 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 464 48 496 792 ;
    LAYER M1 ;
      RECT 464 888 496 1128 ;
    LAYER M1 ;
      RECT 464 1644 496 1884 ;
    LAYER M1 ;
      RECT 544 48 576 792 ;
    LAYER M1 ;
      RECT 624 48 656 792 ;
    LAYER M1 ;
      RECT 624 888 656 1128 ;
    LAYER M1 ;
      RECT 624 1644 656 1884 ;
    LAYER M1 ;
      RECT 704 48 736 792 ;
    LAYER M1 ;
      RECT 784 48 816 792 ;
    LAYER M1 ;
      RECT 784 888 816 1128 ;
    LAYER M1 ;
      RECT 784 1644 816 1884 ;
    LAYER M1 ;
      RECT 864 48 896 792 ;
    LAYER M1 ;
      RECT 944 48 976 792 ;
    LAYER M1 ;
      RECT 944 888 976 1128 ;
    LAYER M1 ;
      RECT 944 1644 976 1884 ;
    LAYER M1 ;
      RECT 1024 48 1056 792 ;
    LAYER M1 ;
      RECT 1104 48 1136 792 ;
    LAYER M1 ;
      RECT 1104 888 1136 1128 ;
    LAYER M1 ;
      RECT 1104 1644 1136 1884 ;
    LAYER M1 ;
      RECT 1184 48 1216 792 ;
    LAYER M2 ;
      RECT 444 68 996 100 ;
    LAYER M2 ;
      RECT 284 908 1156 940 ;
    LAYER M2 ;
      RECT 284 1748 1156 1780 ;
    LAYER M2 ;
      RECT 204 236 1236 268 ;
    LAYER V1 ;
      RECT 624 68 656 100 ;
    LAYER V1 ;
      RECT 624 908 656 940 ;
    LAYER V1 ;
      RECT 624 1748 656 1780 ;
    LAYER V1 ;
      RECT 784 68 816 100 ;
    LAYER V1 ;
      RECT 784 908 816 940 ;
    LAYER V1 ;
      RECT 784 1748 816 1780 ;
    LAYER V1 ;
      RECT 944 68 976 100 ;
    LAYER V1 ;
      RECT 944 908 976 940 ;
    LAYER V1 ;
      RECT 944 1748 976 1780 ;
    LAYER V1 ;
      RECT 464 68 496 100 ;
    LAYER V1 ;
      RECT 464 908 496 940 ;
    LAYER V1 ;
      RECT 464 1748 496 1780 ;
    LAYER V1 ;
      RECT 304 152 336 184 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1748 336 1780 ;
    LAYER V1 ;
      RECT 1104 152 1136 184 ;
    LAYER V1 ;
      RECT 1104 908 1136 940 ;
    LAYER V1 ;
      RECT 1104 1748 1136 1780 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 544 236 576 268 ;
    LAYER V1 ;
      RECT 704 236 736 268 ;
    LAYER V1 ;
      RECT 864 236 896 268 ;
    LAYER V1 ;
      RECT 1024 236 1056 268 ;
    LAYER V1 ;
      RECT 1184 236 1216 268 ;
    LAYER V2 ;
      RECT 464 68 496 100 ;
    LAYER V2 ;
      RECT 464 908 496 940 ;
    LAYER V2 ;
      RECT 624 236 656 268 ;
    LAYER V2 ;
      RECT 624 1748 656 1780 ;
    LAYER V0 ;
      RECT 304 461 336 493 ;
    LAYER V0 ;
      RECT 304 545 336 577 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1748 336 1780 ;
    LAYER V0 ;
      RECT 224 461 256 493 ;
    LAYER V0 ;
      RECT 224 545 256 577 ;
    LAYER V0 ;
      RECT 384 461 416 493 ;
    LAYER V0 ;
      RECT 384 461 416 493 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 464 461 496 493 ;
    LAYER V0 ;
      RECT 464 545 496 577 ;
    LAYER V0 ;
      RECT 464 908 496 940 ;
    LAYER V0 ;
      RECT 464 1748 496 1780 ;
    LAYER V0 ;
      RECT 544 461 576 493 ;
    LAYER V0 ;
      RECT 544 461 576 493 ;
    LAYER V0 ;
      RECT 544 545 576 577 ;
    LAYER V0 ;
      RECT 544 545 576 577 ;
    LAYER V0 ;
      RECT 624 461 656 493 ;
    LAYER V0 ;
      RECT 624 545 656 577 ;
    LAYER V0 ;
      RECT 624 908 656 940 ;
    LAYER V0 ;
      RECT 624 1748 656 1780 ;
    LAYER V0 ;
      RECT 704 461 736 493 ;
    LAYER V0 ;
      RECT 704 461 736 493 ;
    LAYER V0 ;
      RECT 704 545 736 577 ;
    LAYER V0 ;
      RECT 704 545 736 577 ;
    LAYER V0 ;
      RECT 784 461 816 493 ;
    LAYER V0 ;
      RECT 784 545 816 577 ;
    LAYER V0 ;
      RECT 784 908 816 940 ;
    LAYER V0 ;
      RECT 784 1748 816 1780 ;
    LAYER V0 ;
      RECT 864 461 896 493 ;
    LAYER V0 ;
      RECT 864 461 896 493 ;
    LAYER V0 ;
      RECT 864 545 896 577 ;
    LAYER V0 ;
      RECT 864 545 896 577 ;
    LAYER V0 ;
      RECT 944 461 976 493 ;
    LAYER V0 ;
      RECT 944 545 976 577 ;
    LAYER V0 ;
      RECT 944 908 976 940 ;
    LAYER V0 ;
      RECT 944 1748 976 1780 ;
    LAYER V0 ;
      RECT 1024 461 1056 493 ;
    LAYER V0 ;
      RECT 1024 461 1056 493 ;
    LAYER V0 ;
      RECT 1024 545 1056 577 ;
    LAYER V0 ;
      RECT 1024 545 1056 577 ;
    LAYER V0 ;
      RECT 1104 461 1136 493 ;
    LAYER V0 ;
      RECT 1104 545 1136 577 ;
    LAYER V0 ;
      RECT 1104 908 1136 940 ;
    LAYER V0 ;
      RECT 1104 1748 1136 1780 ;
    LAYER V0 ;
      RECT 1184 461 1216 493 ;
    LAYER V0 ;
      RECT 1184 545 1216 577 ;
  END
END SCM_NMOS_57551371
