MACRO TELESCOPIC_OTA_PG0
  ORIGIN 0 0 ;
  FOREIGN TELESCOPIC_OTA_PG0 0 0 ;
  SIZE 1.44 BY 12.936 ;
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 0.46 1.392 0.5 2.304 ;
    END
  END D1
  PIN VBIASP1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.604 6.116 0.836 6.148 ;
    END
  END VBIASP1
  PIN VOUTN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.364 9.308 0.596 9.34 ;
      LAYER M3 ;
        RECT 0.78 9.54 0.82 10.788 ;
      LAYER M2 ;
        RECT 0.56 9.308 0.64 9.34 ;
      LAYER M3 ;
        RECT 0.62 9.219 0.66 9.429 ;
      LAYER M4 ;
        RECT 0.64 9.304 0.8 9.344 ;
      LAYER M3 ;
        RECT 0.78 9.324 0.82 9.576 ;
    END
  END VOUTN
  PIN VOUTP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.844 9.308 1.076 9.34 ;
      LAYER M3 ;
        RECT 0.86 9.456 0.9 10.704 ;
      LAYER M2 ;
        RECT 0.844 9.308 0.916 9.34 ;
      LAYER M3 ;
        RECT 0.86 9.324 0.9 9.492 ;
    END
  END VOUTP
  PIN VBIASP2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.364 8.468 0.596 8.5 ;
      LAYER M2 ;
        RECT 0.844 8.468 1.076 8.5 ;
      LAYER M2 ;
        RECT 0.56 8.468 0.88 8.5 ;
    END
  END VBIASP2
  PIN VBIASN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 0.54 10.296 0.58 11.544 ;
    END
  END VBIASN
  PIN VINP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.444 3.764 1.156 3.796 ;
    END
  END VINP
  PIN VINN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.284 3.68 0.996 3.712 ;
    END
  END VINN
  OBS 
  LAYER M2 ;
        RECT 0.284 2.168 1.156 2.2 ;
  LAYER M2 ;
        RECT 0.204 4.436 1.236 4.468 ;
  LAYER M2 ;
        RECT 0.684 2.168 0.756 2.2 ;
  LAYER M3 ;
        RECT 0.7 2.184 0.74 4.452 ;
  LAYER M2 ;
        RECT 0.684 4.436 0.756 4.468 ;
  LAYER M2 ;
        RECT 0.684 4.436 0.756 4.468 ;
  LAYER M3 ;
        RECT 0.7 4.416 0.74 4.488 ;
  LAYER M2 ;
        RECT 0.684 2.168 0.756 2.2 ;
  LAYER M3 ;
        RECT 0.7 2.148 0.74 2.22 ;
  LAYER M2 ;
        RECT 0.684 4.436 0.756 4.468 ;
  LAYER M3 ;
        RECT 0.7 4.416 0.74 4.488 ;
  LAYER M2 ;
        RECT 0.684 2.168 0.756 2.2 ;
  LAYER M3 ;
        RECT 0.7 2.148 0.74 2.22 ;
  LAYER M2 ;
        RECT 0.444 6.956 0.676 6.988 ;
  LAYER M3 ;
        RECT 0.46 7.608 0.5 9.276 ;
  LAYER M2 ;
        RECT 0.444 6.956 0.516 6.988 ;
  LAYER M3 ;
        RECT 0.46 6.972 0.5 7.644 ;
  LAYER M2 ;
        RECT 0.444 6.956 0.516 6.988 ;
  LAYER M3 ;
        RECT 0.46 6.936 0.5 7.008 ;
  LAYER M2 ;
        RECT 0.444 6.956 0.516 6.988 ;
  LAYER M3 ;
        RECT 0.46 6.936 0.5 7.008 ;
  LAYER M2 ;
        RECT 0.604 6.872 0.836 6.904 ;
  LAYER M3 ;
        RECT 0.94 7.608 0.98 9.276 ;
  LAYER M2 ;
        RECT 0.8 6.872 0.96 6.904 ;
  LAYER M3 ;
        RECT 0.94 6.888 0.98 7.644 ;
  LAYER M2 ;
        RECT 0.924 6.872 0.996 6.904 ;
  LAYER M3 ;
        RECT 0.94 6.852 0.98 6.924 ;
  LAYER M2 ;
        RECT 0.924 6.872 0.996 6.904 ;
  LAYER M3 ;
        RECT 0.94 6.852 0.98 6.924 ;
  LAYER M3 ;
        RECT 0.7 9.624 0.74 10.872 ;
  LAYER M2 ;
        RECT 0.284 4.52 0.996 4.552 ;
  LAYER M3 ;
        RECT 0.7 9.072 0.74 9.66 ;
  LAYER M2 ;
        RECT 0.58 9.056 0.78 9.088 ;
  LAYER M3 ;
        RECT 0.62 4.536 0.66 9.072 ;
  LAYER M2 ;
        RECT 0.604 4.52 0.676 4.552 ;
  LAYER M2 ;
        RECT 0.684 9.056 0.756 9.088 ;
  LAYER M3 ;
        RECT 0.7 9.036 0.74 9.108 ;
  LAYER M2 ;
        RECT 0.604 9.056 0.676 9.088 ;
  LAYER M3 ;
        RECT 0.62 9.036 0.66 9.108 ;
  LAYER M2 ;
        RECT 0.604 4.52 0.676 4.552 ;
  LAYER M3 ;
        RECT 0.62 4.5 0.66 4.572 ;
  LAYER M2 ;
        RECT 0.604 4.52 0.676 4.552 ;
  LAYER M3 ;
        RECT 0.62 4.5 0.66 4.572 ;
  LAYER M3 ;
        RECT 0.62 9.708 0.66 10.956 ;
  LAYER M2 ;
        RECT 0.444 4.604 1.156 4.636 ;
  LAYER M3 ;
        RECT 0.62 9.704 0.66 9.784 ;
  LAYER M4 ;
        RECT 0.53 9.724 0.67 9.764 ;
  LAYER M3 ;
        RECT 0.54 4.62 0.58 9.744 ;
  LAYER M2 ;
        RECT 0.524 4.604 0.596 4.636 ;
  LAYER M2 ;
        RECT 0.524 4.604 0.596 4.636 ;
  LAYER M3 ;
        RECT 0.54 4.584 0.58 4.656 ;
  LAYER M3 ;
        RECT 0.62 9.704 0.66 9.784 ;
  LAYER M4 ;
        RECT 0.6 9.724 0.68 9.764 ;
  LAYER M3 ;
        RECT 0.54 9.704 0.58 9.784 ;
  LAYER M4 ;
        RECT 0.52 9.724 0.6 9.764 ;
  LAYER M2 ;
        RECT 0.524 4.604 0.596 4.636 ;
  LAYER M3 ;
        RECT 0.54 4.584 0.58 4.656 ;
  LAYER M1 ;
        RECT 0.304 1.56 0.336 2.304 ;
  LAYER M1 ;
        RECT 0.304 1.224 0.336 1.464 ;
  LAYER M1 ;
        RECT 0.304 0.468 0.336 0.708 ;
  LAYER M1 ;
        RECT 0.224 1.56 0.256 2.304 ;
  LAYER M1 ;
        RECT 0.384 1.56 0.416 2.304 ;
  LAYER M1 ;
        RECT 0.464 1.56 0.496 2.304 ;
  LAYER M1 ;
        RECT 0.464 1.224 0.496 1.464 ;
  LAYER M1 ;
        RECT 0.464 0.468 0.496 0.708 ;
  LAYER M1 ;
        RECT 0.544 1.56 0.576 2.304 ;
  LAYER M1 ;
        RECT 0.624 1.56 0.656 2.304 ;
  LAYER M1 ;
        RECT 0.624 1.224 0.656 1.464 ;
  LAYER M1 ;
        RECT 0.624 0.468 0.656 0.708 ;
  LAYER M1 ;
        RECT 0.704 1.56 0.736 2.304 ;
  LAYER M1 ;
        RECT 0.784 1.56 0.816 2.304 ;
  LAYER M1 ;
        RECT 0.784 1.224 0.816 1.464 ;
  LAYER M1 ;
        RECT 0.784 0.468 0.816 0.708 ;
  LAYER M1 ;
        RECT 0.864 1.56 0.896 2.304 ;
  LAYER M1 ;
        RECT 0.944 1.56 0.976 2.304 ;
  LAYER M1 ;
        RECT 0.944 1.224 0.976 1.464 ;
  LAYER M1 ;
        RECT 0.944 0.468 0.976 0.708 ;
  LAYER M1 ;
        RECT 1.024 1.56 1.056 2.304 ;
  LAYER M1 ;
        RECT 1.104 1.56 1.136 2.304 ;
  LAYER M1 ;
        RECT 1.104 1.224 1.136 1.464 ;
  LAYER M1 ;
        RECT 1.104 0.468 1.136 0.708 ;
  LAYER M1 ;
        RECT 1.184 1.56 1.216 2.304 ;
  LAYER M2 ;
        RECT 0.444 2.252 0.996 2.284 ;
  LAYER M2 ;
        RECT 0.284 1.412 1.156 1.444 ;
  LAYER M2 ;
        RECT 0.284 0.572 1.156 0.604 ;
  LAYER M2 ;
        RECT 0.204 2.084 1.236 2.116 ;
  LAYER M3 ;
        RECT 0.46 1.392 0.5 2.304 ;
  LAYER M2 ;
        RECT 0.284 2.168 1.156 2.2 ;
  LAYER M3 ;
        RECT 0.62 0.552 0.66 2.136 ;
  LAYER M1 ;
        RECT 0.624 6.264 0.656 7.008 ;
  LAYER M1 ;
        RECT 0.624 5.928 0.656 6.168 ;
  LAYER M1 ;
        RECT 0.624 5.172 0.656 5.412 ;
  LAYER M1 ;
        RECT 0.544 6.264 0.576 7.008 ;
  LAYER M1 ;
        RECT 0.704 6.264 0.736 7.008 ;
  LAYER M1 ;
        RECT 0.784 6.264 0.816 7.008 ;
  LAYER M1 ;
        RECT 0.784 5.928 0.816 6.168 ;
  LAYER M1 ;
        RECT 0.784 5.172 0.816 5.412 ;
  LAYER M1 ;
        RECT 0.864 6.264 0.896 7.008 ;
  LAYER M2 ;
        RECT 0.604 5.276 0.836 5.308 ;
  LAYER M2 ;
        RECT 0.524 6.788 0.916 6.82 ;
  LAYER M2 ;
        RECT 0.444 6.956 0.676 6.988 ;
  LAYER M2 ;
        RECT 0.604 6.872 0.836 6.904 ;
  LAYER M2 ;
        RECT 0.604 6.116 0.836 6.148 ;
  LAYER M3 ;
        RECT 0.7 5.256 0.74 6.84 ;
  LAYER M1 ;
        RECT 0.384 8.616 0.416 9.36 ;
  LAYER M1 ;
        RECT 0.384 8.28 0.416 8.52 ;
  LAYER M1 ;
        RECT 0.384 7.524 0.416 7.764 ;
  LAYER M1 ;
        RECT 0.464 8.616 0.496 9.36 ;
  LAYER M1 ;
        RECT 0.304 8.616 0.336 9.36 ;
  LAYER M2 ;
        RECT 0.364 7.628 0.596 7.66 ;
  LAYER M2 ;
        RECT 0.284 9.224 0.516 9.256 ;
  LAYER M2 ;
        RECT 0.364 9.308 0.596 9.34 ;
  LAYER M2 ;
        RECT 0.364 8.468 0.596 8.5 ;
  LAYER M3 ;
        RECT 0.46 7.608 0.5 9.276 ;
  LAYER M1 ;
        RECT 1.024 8.616 1.056 9.36 ;
  LAYER M1 ;
        RECT 1.024 8.28 1.056 8.52 ;
  LAYER M1 ;
        RECT 1.024 7.524 1.056 7.764 ;
  LAYER M1 ;
        RECT 0.944 8.616 0.976 9.36 ;
  LAYER M1 ;
        RECT 1.104 8.616 1.136 9.36 ;
  LAYER M2 ;
        RECT 0.844 7.628 1.076 7.66 ;
  LAYER M2 ;
        RECT 0.924 9.224 1.156 9.256 ;
  LAYER M2 ;
        RECT 0.844 9.308 1.076 9.34 ;
  LAYER M2 ;
        RECT 0.844 8.468 1.076 8.5 ;
  LAYER M3 ;
        RECT 0.94 7.608 0.98 9.276 ;
  LAYER M1 ;
        RECT 1.024 9.456 1.056 10.2 ;
  LAYER M1 ;
        RECT 1.024 10.296 1.056 10.536 ;
  LAYER M1 ;
        RECT 1.024 10.632 1.056 11.376 ;
  LAYER M1 ;
        RECT 1.024 11.472 1.056 11.712 ;
  LAYER M1 ;
        RECT 1.024 12.228 1.056 12.468 ;
  LAYER M1 ;
        RECT 1.104 9.456 1.136 10.2 ;
  LAYER M1 ;
        RECT 1.104 10.632 1.136 11.376 ;
  LAYER M1 ;
        RECT 0.944 9.456 0.976 10.2 ;
  LAYER M1 ;
        RECT 0.944 10.632 0.976 11.376 ;
  LAYER M1 ;
        RECT 0.384 9.456 0.416 10.2 ;
  LAYER M1 ;
        RECT 0.384 10.296 0.416 10.536 ;
  LAYER M1 ;
        RECT 0.384 10.632 0.416 11.376 ;
  LAYER M1 ;
        RECT 0.384 11.472 0.416 11.712 ;
  LAYER M1 ;
        RECT 0.384 12.228 0.416 12.468 ;
  LAYER M1 ;
        RECT 0.464 9.456 0.496 10.2 ;
  LAYER M1 ;
        RECT 0.464 10.632 0.496 11.376 ;
  LAYER M1 ;
        RECT 0.304 9.456 0.336 10.2 ;
  LAYER M1 ;
        RECT 0.304 10.632 0.336 11.376 ;
  LAYER M2 ;
        RECT 0.844 9.476 1.076 9.508 ;
  LAYER M2 ;
        RECT 0.364 9.56 0.836 9.592 ;
  LAYER M2 ;
        RECT 0.684 9.644 1.156 9.676 ;
  LAYER M2 ;
        RECT 0.284 9.728 0.676 9.76 ;
  LAYER M2 ;
        RECT 0.364 10.316 1.076 10.348 ;
  LAYER M2 ;
        RECT 0.364 10.652 0.916 10.684 ;
  LAYER M2 ;
        RECT 0.764 10.736 1.076 10.768 ;
  LAYER M2 ;
        RECT 0.284 10.82 0.756 10.852 ;
  LAYER M2 ;
        RECT 0.604 10.904 1.156 10.936 ;
  LAYER M2 ;
        RECT 0.364 11.492 1.076 11.524 ;
  LAYER M2 ;
        RECT 0.364 12.332 1.076 12.364 ;
  LAYER M3 ;
        RECT 0.86 9.456 0.9 10.704 ;
  LAYER M3 ;
        RECT 0.78 9.54 0.82 10.788 ;
  LAYER M3 ;
        RECT 0.54 10.296 0.58 11.544 ;
  LAYER M3 ;
        RECT 0.7 9.624 0.74 10.872 ;
  LAYER M3 ;
        RECT 0.62 9.708 0.66 10.956 ;
  LAYER M1 ;
        RECT 1.104 3.912 1.136 4.656 ;
  LAYER M1 ;
        RECT 1.104 3.576 1.136 3.816 ;
  LAYER M1 ;
        RECT 1.104 2.82 1.136 3.06 ;
  LAYER M1 ;
        RECT 1.184 3.912 1.216 4.656 ;
  LAYER M1 ;
        RECT 1.024 3.912 1.056 4.656 ;
  LAYER M1 ;
        RECT 0.944 3.912 0.976 4.656 ;
  LAYER M1 ;
        RECT 0.944 3.576 0.976 3.816 ;
  LAYER M1 ;
        RECT 0.944 2.82 0.976 3.06 ;
  LAYER M1 ;
        RECT 0.864 3.912 0.896 4.656 ;
  LAYER M1 ;
        RECT 0.784 3.912 0.816 4.656 ;
  LAYER M1 ;
        RECT 0.784 3.576 0.816 3.816 ;
  LAYER M1 ;
        RECT 0.784 2.82 0.816 3.06 ;
  LAYER M1 ;
        RECT 0.704 3.912 0.736 4.656 ;
  LAYER M1 ;
        RECT 0.624 3.912 0.656 4.656 ;
  LAYER M1 ;
        RECT 0.624 3.576 0.656 3.816 ;
  LAYER M1 ;
        RECT 0.624 2.82 0.656 3.06 ;
  LAYER M1 ;
        RECT 0.544 3.912 0.576 4.656 ;
  LAYER M1 ;
        RECT 0.464 3.912 0.496 4.656 ;
  LAYER M1 ;
        RECT 0.464 3.576 0.496 3.816 ;
  LAYER M1 ;
        RECT 0.464 2.82 0.496 3.06 ;
  LAYER M1 ;
        RECT 0.384 3.912 0.416 4.656 ;
  LAYER M1 ;
        RECT 0.304 3.912 0.336 4.656 ;
  LAYER M1 ;
        RECT 0.304 3.576 0.336 3.816 ;
  LAYER M1 ;
        RECT 0.304 2.82 0.336 3.06 ;
  LAYER M1 ;
        RECT 0.224 3.912 0.256 4.656 ;
  LAYER M2 ;
        RECT 0.284 2.924 1.156 2.956 ;
  LAYER M2 ;
        RECT 0.444 4.604 1.156 4.636 ;
  LAYER M2 ;
        RECT 0.284 4.52 0.996 4.552 ;
  LAYER M2 ;
        RECT 0.444 3.764 1.156 3.796 ;
  LAYER M2 ;
        RECT 0.284 3.68 0.996 3.712 ;
  LAYER M2 ;
        RECT 0.204 4.436 1.236 4.468 ;
  END 
END TELESCOPIC_OTA_PG0
