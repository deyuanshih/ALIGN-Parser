MACRO SCM_NMOS_57551371
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_57551371 0 0 ;
  SIZE 1440 BY 2352 ;
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 460 48 500 960 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 152 1156 184 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 620 216 660 1800 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1644 336 1884 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 464 48 496 792 ;
    LAYER M1 ;
      RECT 464 888 496 1128 ;
    LAYER M1 ;
      RECT 464 1644 496 1884 ;
    LAYER M1 ;
      RECT 544 48 576 792 ;
    LAYER M1 ;
      RECT 624 48 656 792 ;
    LAYER M1 ;
      RECT 624 888 656 1128 ;
    LAYER M1 ;
      RECT 624 1644 656 1884 ;
    LAYER M1 ;
      RECT 704 48 736 792 ;
    LAYER M1 ;
      RECT 784 48 816 792 ;
    LAYER M1 ;
      RECT 784 888 816 1128 ;
    LAYER M1 ;
      RECT 784 1644 816 1884 ;
    LAYER M1 ;
      RECT 864 48 896 792 ;
    LAYER M1 ;
      RECT 944 48 976 792 ;
    LAYER M1 ;
      RECT 944 888 976 1128 ;
    LAYER M1 ;
      RECT 944 1644 976 1884 ;
    LAYER M1 ;
      RECT 1024 48 1056 792 ;
    LAYER M1 ;
      RECT 1104 48 1136 792 ;
    LAYER M1 ;
      RECT 1104 888 1136 1128 ;
    LAYER M1 ;
      RECT 1104 1644 1136 1884 ;
    LAYER M1 ;
      RECT 1184 48 1216 792 ;
    LAYER M2 ;
      RECT 444 68 996 100 ;
    LAYER M2 ;
      RECT 284 908 1156 940 ;
    LAYER M2 ;
      RECT 284 1748 1156 1780 ;
    LAYER M2 ;
      RECT 204 236 1236 268 ;
    LAYER V1 ;
      RECT 624 68 656 100 ;
    LAYER V1 ;
      RECT 624 908 656 940 ;
    LAYER V1 ;
      RECT 624 1748 656 1780 ;
    LAYER V1 ;
      RECT 784 68 816 100 ;
    LAYER V1 ;
      RECT 784 908 816 940 ;
    LAYER V1 ;
      RECT 784 1748 816 1780 ;
    LAYER V1 ;
      RECT 944 68 976 100 ;
    LAYER V1 ;
      RECT 944 908 976 940 ;
    LAYER V1 ;
      RECT 944 1748 976 1780 ;
    LAYER V1 ;
      RECT 464 68 496 100 ;
    LAYER V1 ;
      RECT 464 908 496 940 ;
    LAYER V1 ;
      RECT 464 1748 496 1780 ;
    LAYER V1 ;
      RECT 304 152 336 184 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1748 336 1780 ;
    LAYER V1 ;
      RECT 1104 152 1136 184 ;
    LAYER V1 ;
      RECT 1104 908 1136 940 ;
    LAYER V1 ;
      RECT 1104 1748 1136 1780 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 544 236 576 268 ;
    LAYER V1 ;
      RECT 704 236 736 268 ;
    LAYER V1 ;
      RECT 864 236 896 268 ;
    LAYER V1 ;
      RECT 1024 236 1056 268 ;
    LAYER V1 ;
      RECT 1184 236 1216 268 ;
    LAYER V2 ;
      RECT 464 68 496 100 ;
    LAYER V2 ;
      RECT 464 908 496 940 ;
    LAYER V2 ;
      RECT 624 236 656 268 ;
    LAYER V2 ;
      RECT 624 1748 656 1780 ;
    LAYER V0 ;
      RECT 304 461 336 493 ;
    LAYER V0 ;
      RECT 304 545 336 577 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1748 336 1780 ;
    LAYER V0 ;
      RECT 224 461 256 493 ;
    LAYER V0 ;
      RECT 224 545 256 577 ;
    LAYER V0 ;
      RECT 384 461 416 493 ;
    LAYER V0 ;
      RECT 384 461 416 493 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 464 461 496 493 ;
    LAYER V0 ;
      RECT 464 545 496 577 ;
    LAYER V0 ;
      RECT 464 908 496 940 ;
    LAYER V0 ;
      RECT 464 1748 496 1780 ;
    LAYER V0 ;
      RECT 544 461 576 493 ;
    LAYER V0 ;
      RECT 544 461 576 493 ;
    LAYER V0 ;
      RECT 544 545 576 577 ;
    LAYER V0 ;
      RECT 544 545 576 577 ;
    LAYER V0 ;
      RECT 624 461 656 493 ;
    LAYER V0 ;
      RECT 624 545 656 577 ;
    LAYER V0 ;
      RECT 624 908 656 940 ;
    LAYER V0 ;
      RECT 624 1748 656 1780 ;
    LAYER V0 ;
      RECT 704 461 736 493 ;
    LAYER V0 ;
      RECT 704 461 736 493 ;
    LAYER V0 ;
      RECT 704 545 736 577 ;
    LAYER V0 ;
      RECT 704 545 736 577 ;
    LAYER V0 ;
      RECT 784 461 816 493 ;
    LAYER V0 ;
      RECT 784 545 816 577 ;
    LAYER V0 ;
      RECT 784 908 816 940 ;
    LAYER V0 ;
      RECT 784 1748 816 1780 ;
    LAYER V0 ;
      RECT 864 461 896 493 ;
    LAYER V0 ;
      RECT 864 461 896 493 ;
    LAYER V0 ;
      RECT 864 545 896 577 ;
    LAYER V0 ;
      RECT 864 545 896 577 ;
    LAYER V0 ;
      RECT 944 461 976 493 ;
    LAYER V0 ;
      RECT 944 545 976 577 ;
    LAYER V0 ;
      RECT 944 908 976 940 ;
    LAYER V0 ;
      RECT 944 1748 976 1780 ;
    LAYER V0 ;
      RECT 1024 461 1056 493 ;
    LAYER V0 ;
      RECT 1024 461 1056 493 ;
    LAYER V0 ;
      RECT 1024 545 1056 577 ;
    LAYER V0 ;
      RECT 1024 545 1056 577 ;
    LAYER V0 ;
      RECT 1104 461 1136 493 ;
    LAYER V0 ;
      RECT 1104 545 1136 577 ;
    LAYER V0 ;
      RECT 1104 908 1136 940 ;
    LAYER V0 ;
      RECT 1104 1748 1136 1780 ;
    LAYER V0 ;
      RECT 1184 461 1216 493 ;
    LAYER V0 ;
      RECT 1184 545 1216 577 ;
  END
END SCM_NMOS_57551371
MACRO CMC_PMOS_95878848_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_95878848_X1_Y1 0 0 ;
  SIZE 800 BY 2352 ;
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124 68 356 100 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 152 516 184 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 908 516 940 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 380 216 420 1800 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1644 336 1884 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 464 48 496 792 ;
    LAYER M1 ;
      RECT 464 888 496 1128 ;
    LAYER M1 ;
      RECT 464 1644 496 1884 ;
    LAYER M1 ;
      RECT 544 48 576 792 ;
    LAYER M2 ;
      RECT 284 1748 516 1780 ;
    LAYER M2 ;
      RECT 204 236 596 268 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1748 336 1780 ;
    LAYER V1 ;
      RECT 464 152 496 184 ;
    LAYER V1 ;
      RECT 464 908 496 940 ;
    LAYER V1 ;
      RECT 464 1748 496 1780 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 544 236 576 268 ;
    LAYER V2 ;
      RECT 384 236 416 268 ;
    LAYER V2 ;
      RECT 384 1748 416 1780 ;
    LAYER V0 ;
      RECT 304 461 336 493 ;
    LAYER V0 ;
      RECT 304 545 336 577 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1748 336 1780 ;
    LAYER V0 ;
      RECT 224 461 256 493 ;
    LAYER V0 ;
      RECT 224 545 256 577 ;
    LAYER V0 ;
      RECT 384 461 416 493 ;
    LAYER V0 ;
      RECT 384 461 416 493 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 464 461 496 493 ;
    LAYER V0 ;
      RECT 464 545 496 577 ;
    LAYER V0 ;
      RECT 464 908 496 940 ;
    LAYER V0 ;
      RECT 464 1748 496 1780 ;
    LAYER V0 ;
      RECT 544 461 576 493 ;
    LAYER V0 ;
      RECT 544 545 576 577 ;
  END
END CMC_PMOS_95878848_X1_Y1
MACRO CMC_S_NMOS_B_2722902_X1_Y2
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CMC_S_NMOS_B_2722902_X1_Y2 0 0 ;
  SIZE 1280 BY 3528 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 2924 996 2956 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 460 48 500 1296 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 540 132 580 1380 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 780 888 820 2136 ;
    END
  END G
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 620 216 660 1464 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 700 300 740 1548 ;
    END
  END SB
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1224 336 1968 ;
    LAYER M1 ;
      RECT 304 2064 336 2304 ;
    LAYER M1 ;
      RECT 304 2820 336 3060 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 224 1224 256 1968 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 384 1224 416 1968 ;
    LAYER M1 ;
      RECT 944 48 976 792 ;
    LAYER M1 ;
      RECT 944 888 976 1128 ;
    LAYER M1 ;
      RECT 944 1224 976 1968 ;
    LAYER M1 ;
      RECT 944 2064 976 2304 ;
    LAYER M1 ;
      RECT 944 2820 976 3060 ;
    LAYER M1 ;
      RECT 864 48 896 792 ;
    LAYER M1 ;
      RECT 864 1224 896 1968 ;
    LAYER M1 ;
      RECT 1024 48 1056 792 ;
    LAYER M1 ;
      RECT 1024 1224 1056 1968 ;
    LAYER M2 ;
      RECT 284 68 516 100 ;
    LAYER M2 ;
      RECT 524 152 996 184 ;
    LAYER M2 ;
      RECT 204 236 676 268 ;
    LAYER M2 ;
      RECT 684 320 1076 352 ;
    LAYER M2 ;
      RECT 284 908 996 940 ;
    LAYER M2 ;
      RECT 444 1244 996 1276 ;
    LAYER M2 ;
      RECT 284 1328 596 1360 ;
    LAYER M2 ;
      RECT 604 1412 1076 1444 ;
    LAYER M2 ;
      RECT 204 1496 756 1528 ;
    LAYER M2 ;
      RECT 284 2084 996 2116 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1328 336 1360 ;
    LAYER V1 ;
      RECT 304 2084 336 2116 ;
    LAYER V1 ;
      RECT 304 2924 336 2956 ;
    LAYER V1 ;
      RECT 944 152 976 184 ;
    LAYER V1 ;
      RECT 944 908 976 940 ;
    LAYER V1 ;
      RECT 944 1244 976 1276 ;
    LAYER V1 ;
      RECT 944 2084 976 2116 ;
    LAYER V1 ;
      RECT 944 2924 976 2956 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 224 1496 256 1528 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 384 1496 416 1528 ;
    LAYER V1 ;
      RECT 864 320 896 352 ;
    LAYER V1 ;
      RECT 864 1412 896 1444 ;
    LAYER V1 ;
      RECT 1024 320 1056 352 ;
    LAYER V1 ;
      RECT 1024 1412 1056 1444 ;
    LAYER V2 ;
      RECT 464 68 496 100 ;
    LAYER V2 ;
      RECT 464 1244 496 1276 ;
    LAYER V2 ;
      RECT 544 152 576 184 ;
    LAYER V2 ;
      RECT 544 1328 576 1360 ;
    LAYER V2 ;
      RECT 624 236 656 268 ;
    LAYER V2 ;
      RECT 624 1412 656 1444 ;
    LAYER V2 ;
      RECT 704 320 736 352 ;
    LAYER V2 ;
      RECT 704 1496 736 1528 ;
    LAYER V2 ;
      RECT 784 908 816 940 ;
    LAYER V2 ;
      RECT 784 2084 816 2116 ;
    LAYER V0 ;
      RECT 304 398 336 430 ;
    LAYER V0 ;
      RECT 304 482 336 514 ;
    LAYER V0 ;
      RECT 304 566 336 598 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1574 336 1606 ;
    LAYER V0 ;
      RECT 304 1658 336 1690 ;
    LAYER V0 ;
      RECT 304 1742 336 1774 ;
    LAYER V0 ;
      RECT 304 2084 336 2116 ;
    LAYER V0 ;
      RECT 304 2924 336 2956 ;
    LAYER V0 ;
      RECT 304 2924 336 2956 ;
    LAYER V0 ;
      RECT 224 398 256 430 ;
    LAYER V0 ;
      RECT 224 482 256 514 ;
    LAYER V0 ;
      RECT 224 566 256 598 ;
    LAYER V0 ;
      RECT 224 1574 256 1606 ;
    LAYER V0 ;
      RECT 224 1658 256 1690 ;
    LAYER V0 ;
      RECT 224 1742 256 1774 ;
    LAYER V0 ;
      RECT 384 398 416 430 ;
    LAYER V0 ;
      RECT 384 482 416 514 ;
    LAYER V0 ;
      RECT 384 566 416 598 ;
    LAYER V0 ;
      RECT 384 1574 416 1606 ;
    LAYER V0 ;
      RECT 384 1658 416 1690 ;
    LAYER V0 ;
      RECT 384 1742 416 1774 ;
    LAYER V0 ;
      RECT 944 398 976 430 ;
    LAYER V0 ;
      RECT 944 482 976 514 ;
    LAYER V0 ;
      RECT 944 566 976 598 ;
    LAYER V0 ;
      RECT 944 908 976 940 ;
    LAYER V0 ;
      RECT 944 1574 976 1606 ;
    LAYER V0 ;
      RECT 944 1658 976 1690 ;
    LAYER V0 ;
      RECT 944 1742 976 1774 ;
    LAYER V0 ;
      RECT 944 2084 976 2116 ;
    LAYER V0 ;
      RECT 944 2924 976 2956 ;
    LAYER V0 ;
      RECT 944 2924 976 2956 ;
    LAYER V0 ;
      RECT 864 398 896 430 ;
    LAYER V0 ;
      RECT 864 482 896 514 ;
    LAYER V0 ;
      RECT 864 566 896 598 ;
    LAYER V0 ;
      RECT 864 1574 896 1606 ;
    LAYER V0 ;
      RECT 864 1658 896 1690 ;
    LAYER V0 ;
      RECT 864 1742 896 1774 ;
    LAYER V0 ;
      RECT 1024 398 1056 430 ;
    LAYER V0 ;
      RECT 1024 482 1056 514 ;
    LAYER V0 ;
      RECT 1024 566 1056 598 ;
    LAYER V0 ;
      RECT 1024 1574 1056 1606 ;
    LAYER V0 ;
      RECT 1024 1658 1056 1690 ;
    LAYER V0 ;
      RECT 1024 1742 1056 1774 ;
  END
END CMC_S_NMOS_B_2722902_X1_Y2
MACRO CMC_S_NMOS_B_2722902_X2_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CMC_S_NMOS_B_2722902_X2_Y1 0 0 ;
  SIZE 2560 BY 2352 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 1748 2276 1780 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 68 996 100 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1564 152 2276 184 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 908 2276 940 ;
    END
  END G
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204 236 1076 268 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1484 320 2356 352 ;
    END
  END SB
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1644 336 1884 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 944 48 976 792 ;
    LAYER M1 ;
      RECT 944 888 976 1128 ;
    LAYER M1 ;
      RECT 944 1644 976 1884 ;
    LAYER M1 ;
      RECT 864 48 896 792 ;
    LAYER M1 ;
      RECT 1024 48 1056 792 ;
    LAYER M1 ;
      RECT 1584 48 1616 792 ;
    LAYER M1 ;
      RECT 1584 888 1616 1128 ;
    LAYER M1 ;
      RECT 1584 1644 1616 1884 ;
    LAYER M1 ;
      RECT 1504 48 1536 792 ;
    LAYER M1 ;
      RECT 1664 48 1696 792 ;
    LAYER M1 ;
      RECT 2224 48 2256 792 ;
    LAYER M1 ;
      RECT 2224 888 2256 1128 ;
    LAYER M1 ;
      RECT 2224 1644 2256 1884 ;
    LAYER M1 ;
      RECT 2144 48 2176 792 ;
    LAYER M1 ;
      RECT 2304 48 2336 792 ;
    LAYER V1 ;
      RECT 944 68 976 100 ;
    LAYER V1 ;
      RECT 944 908 976 940 ;
    LAYER V1 ;
      RECT 944 1748 976 1780 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1748 336 1780 ;
    LAYER V1 ;
      RECT 2224 152 2256 184 ;
    LAYER V1 ;
      RECT 2224 908 2256 940 ;
    LAYER V1 ;
      RECT 2224 1748 2256 1780 ;
    LAYER V1 ;
      RECT 1584 152 1616 184 ;
    LAYER V1 ;
      RECT 1584 908 1616 940 ;
    LAYER V1 ;
      RECT 1584 1748 1616 1780 ;
    LAYER V1 ;
      RECT 864 236 896 268 ;
    LAYER V1 ;
      RECT 1024 236 1056 268 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 2144 320 2176 352 ;
    LAYER V1 ;
      RECT 1664 320 1696 352 ;
    LAYER V1 ;
      RECT 1504 320 1536 352 ;
    LAYER V1 ;
      RECT 2304 320 2336 352 ;
    LAYER V0 ;
      RECT 304 398 336 430 ;
    LAYER V0 ;
      RECT 304 482 336 514 ;
    LAYER V0 ;
      RECT 304 566 336 598 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1748 336 1780 ;
    LAYER V0 ;
      RECT 224 398 256 430 ;
    LAYER V0 ;
      RECT 224 482 256 514 ;
    LAYER V0 ;
      RECT 224 566 256 598 ;
    LAYER V0 ;
      RECT 384 398 416 430 ;
    LAYER V0 ;
      RECT 384 482 416 514 ;
    LAYER V0 ;
      RECT 384 566 416 598 ;
    LAYER V0 ;
      RECT 944 398 976 430 ;
    LAYER V0 ;
      RECT 944 482 976 514 ;
    LAYER V0 ;
      RECT 944 566 976 598 ;
    LAYER V0 ;
      RECT 944 908 976 940 ;
    LAYER V0 ;
      RECT 944 1748 976 1780 ;
    LAYER V0 ;
      RECT 864 398 896 430 ;
    LAYER V0 ;
      RECT 864 482 896 514 ;
    LAYER V0 ;
      RECT 864 566 896 598 ;
    LAYER V0 ;
      RECT 1024 398 1056 430 ;
    LAYER V0 ;
      RECT 1024 482 1056 514 ;
    LAYER V0 ;
      RECT 1024 566 1056 598 ;
    LAYER V0 ;
      RECT 1584 398 1616 430 ;
    LAYER V0 ;
      RECT 1584 482 1616 514 ;
    LAYER V0 ;
      RECT 1584 566 1616 598 ;
    LAYER V0 ;
      RECT 1584 908 1616 940 ;
    LAYER V0 ;
      RECT 1584 1748 1616 1780 ;
    LAYER V0 ;
      RECT 1504 398 1536 430 ;
    LAYER V0 ;
      RECT 1504 482 1536 514 ;
    LAYER V0 ;
      RECT 1504 566 1536 598 ;
    LAYER V0 ;
      RECT 1664 398 1696 430 ;
    LAYER V0 ;
      RECT 1664 482 1696 514 ;
    LAYER V0 ;
      RECT 1664 566 1696 598 ;
    LAYER V0 ;
      RECT 2224 398 2256 430 ;
    LAYER V0 ;
      RECT 2224 482 2256 514 ;
    LAYER V0 ;
      RECT 2224 566 2256 598 ;
    LAYER V0 ;
      RECT 2224 908 2256 940 ;
    LAYER V0 ;
      RECT 2224 1748 2256 1780 ;
    LAYER V0 ;
      RECT 2144 398 2176 430 ;
    LAYER V0 ;
      RECT 2144 482 2176 514 ;
    LAYER V0 ;
      RECT 2144 566 2176 598 ;
    LAYER V0 ;
      RECT 2304 398 2336 430 ;
    LAYER V0 ;
      RECT 2304 482 2336 514 ;
    LAYER V0 ;
      RECT 2304 566 2336 598 ;
  END
END CMC_S_NMOS_B_2722902_X2_Y1
MACRO DP_NMOS_B_40344802_X3_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_40344802_X3_Y1 0 0 ;
  SIZE 1440 BY 2352 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 1748 1156 1780 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 68 996 100 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 444 152 1156 184 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 908 996 940 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 444 992 1156 1024 ;
    END
  END GB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204 236 1236 268 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1644 336 1884 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 464 48 496 792 ;
    LAYER M1 ;
      RECT 464 888 496 1128 ;
    LAYER M1 ;
      RECT 464 1644 496 1884 ;
    LAYER M1 ;
      RECT 544 48 576 792 ;
    LAYER M1 ;
      RECT 624 48 656 792 ;
    LAYER M1 ;
      RECT 624 888 656 1128 ;
    LAYER M1 ;
      RECT 624 1644 656 1884 ;
    LAYER M1 ;
      RECT 704 48 736 792 ;
    LAYER M1 ;
      RECT 784 48 816 792 ;
    LAYER M1 ;
      RECT 784 888 816 1128 ;
    LAYER M1 ;
      RECT 784 1644 816 1884 ;
    LAYER M1 ;
      RECT 864 48 896 792 ;
    LAYER M1 ;
      RECT 944 48 976 792 ;
    LAYER M1 ;
      RECT 944 888 976 1128 ;
    LAYER M1 ;
      RECT 944 1644 976 1884 ;
    LAYER M1 ;
      RECT 1024 48 1056 792 ;
    LAYER M1 ;
      RECT 1104 48 1136 792 ;
    LAYER M1 ;
      RECT 1104 888 1136 1128 ;
    LAYER M1 ;
      RECT 1104 1644 1136 1884 ;
    LAYER M1 ;
      RECT 1184 48 1216 792 ;
    LAYER V1 ;
      RECT 624 68 656 100 ;
    LAYER V1 ;
      RECT 624 908 656 940 ;
    LAYER V1 ;
      RECT 624 1748 656 1780 ;
    LAYER V1 ;
      RECT 944 68 976 100 ;
    LAYER V1 ;
      RECT 944 908 976 940 ;
    LAYER V1 ;
      RECT 944 1748 976 1780 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1748 336 1780 ;
    LAYER V1 ;
      RECT 784 152 816 184 ;
    LAYER V1 ;
      RECT 784 992 816 1024 ;
    LAYER V1 ;
      RECT 784 1748 816 1780 ;
    LAYER V1 ;
      RECT 464 152 496 184 ;
    LAYER V1 ;
      RECT 464 992 496 1024 ;
    LAYER V1 ;
      RECT 464 1748 496 1780 ;
    LAYER V1 ;
      RECT 1104 152 1136 184 ;
    LAYER V1 ;
      RECT 1104 992 1136 1024 ;
    LAYER V1 ;
      RECT 1104 1748 1136 1780 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 544 236 576 268 ;
    LAYER V1 ;
      RECT 704 236 736 268 ;
    LAYER V1 ;
      RECT 864 236 896 268 ;
    LAYER V1 ;
      RECT 1024 236 1056 268 ;
    LAYER V1 ;
      RECT 1184 236 1216 268 ;
    LAYER V0 ;
      RECT 304 335 336 367 ;
    LAYER V0 ;
      RECT 304 419 336 451 ;
    LAYER V0 ;
      RECT 304 503 336 535 ;
    LAYER V0 ;
      RECT 304 587 336 619 ;
    LAYER V0 ;
      RECT 304 671 336 703 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1748 336 1780 ;
    LAYER V0 ;
      RECT 224 335 256 367 ;
    LAYER V0 ;
      RECT 224 419 256 451 ;
    LAYER V0 ;
      RECT 224 503 256 535 ;
    LAYER V0 ;
      RECT 224 587 256 619 ;
    LAYER V0 ;
      RECT 224 671 256 703 ;
    LAYER V0 ;
      RECT 384 335 416 367 ;
    LAYER V0 ;
      RECT 384 335 416 367 ;
    LAYER V0 ;
      RECT 384 419 416 451 ;
    LAYER V0 ;
      RECT 384 419 416 451 ;
    LAYER V0 ;
      RECT 384 503 416 535 ;
    LAYER V0 ;
      RECT 384 503 416 535 ;
    LAYER V0 ;
      RECT 384 587 416 619 ;
    LAYER V0 ;
      RECT 384 587 416 619 ;
    LAYER V0 ;
      RECT 384 671 416 703 ;
    LAYER V0 ;
      RECT 384 671 416 703 ;
    LAYER V0 ;
      RECT 464 335 496 367 ;
    LAYER V0 ;
      RECT 464 419 496 451 ;
    LAYER V0 ;
      RECT 464 503 496 535 ;
    LAYER V0 ;
      RECT 464 587 496 619 ;
    LAYER V0 ;
      RECT 464 671 496 703 ;
    LAYER V0 ;
      RECT 464 908 496 940 ;
    LAYER V0 ;
      RECT 464 1748 496 1780 ;
    LAYER V0 ;
      RECT 544 335 576 367 ;
    LAYER V0 ;
      RECT 544 335 576 367 ;
    LAYER V0 ;
      RECT 544 419 576 451 ;
    LAYER V0 ;
      RECT 544 419 576 451 ;
    LAYER V0 ;
      RECT 544 503 576 535 ;
    LAYER V0 ;
      RECT 544 503 576 535 ;
    LAYER V0 ;
      RECT 544 587 576 619 ;
    LAYER V0 ;
      RECT 544 587 576 619 ;
    LAYER V0 ;
      RECT 544 671 576 703 ;
    LAYER V0 ;
      RECT 544 671 576 703 ;
    LAYER V0 ;
      RECT 624 335 656 367 ;
    LAYER V0 ;
      RECT 624 419 656 451 ;
    LAYER V0 ;
      RECT 624 503 656 535 ;
    LAYER V0 ;
      RECT 624 587 656 619 ;
    LAYER V0 ;
      RECT 624 671 656 703 ;
    LAYER V0 ;
      RECT 624 908 656 940 ;
    LAYER V0 ;
      RECT 624 1748 656 1780 ;
    LAYER V0 ;
      RECT 704 335 736 367 ;
    LAYER V0 ;
      RECT 704 335 736 367 ;
    LAYER V0 ;
      RECT 704 419 736 451 ;
    LAYER V0 ;
      RECT 704 419 736 451 ;
    LAYER V0 ;
      RECT 704 503 736 535 ;
    LAYER V0 ;
      RECT 704 503 736 535 ;
    LAYER V0 ;
      RECT 704 587 736 619 ;
    LAYER V0 ;
      RECT 704 587 736 619 ;
    LAYER V0 ;
      RECT 704 671 736 703 ;
    LAYER V0 ;
      RECT 704 671 736 703 ;
    LAYER V0 ;
      RECT 784 335 816 367 ;
    LAYER V0 ;
      RECT 784 419 816 451 ;
    LAYER V0 ;
      RECT 784 503 816 535 ;
    LAYER V0 ;
      RECT 784 587 816 619 ;
    LAYER V0 ;
      RECT 784 671 816 703 ;
    LAYER V0 ;
      RECT 784 908 816 940 ;
    LAYER V0 ;
      RECT 784 1748 816 1780 ;
    LAYER V0 ;
      RECT 864 335 896 367 ;
    LAYER V0 ;
      RECT 864 335 896 367 ;
    LAYER V0 ;
      RECT 864 419 896 451 ;
    LAYER V0 ;
      RECT 864 419 896 451 ;
    LAYER V0 ;
      RECT 864 503 896 535 ;
    LAYER V0 ;
      RECT 864 503 896 535 ;
    LAYER V0 ;
      RECT 864 587 896 619 ;
    LAYER V0 ;
      RECT 864 587 896 619 ;
    LAYER V0 ;
      RECT 864 671 896 703 ;
    LAYER V0 ;
      RECT 864 671 896 703 ;
    LAYER V0 ;
      RECT 944 335 976 367 ;
    LAYER V0 ;
      RECT 944 419 976 451 ;
    LAYER V0 ;
      RECT 944 503 976 535 ;
    LAYER V0 ;
      RECT 944 587 976 619 ;
    LAYER V0 ;
      RECT 944 671 976 703 ;
    LAYER V0 ;
      RECT 944 908 976 940 ;
    LAYER V0 ;
      RECT 944 1748 976 1780 ;
    LAYER V0 ;
      RECT 1024 335 1056 367 ;
    LAYER V0 ;
      RECT 1024 335 1056 367 ;
    LAYER V0 ;
      RECT 1024 419 1056 451 ;
    LAYER V0 ;
      RECT 1024 419 1056 451 ;
    LAYER V0 ;
      RECT 1024 503 1056 535 ;
    LAYER V0 ;
      RECT 1024 503 1056 535 ;
    LAYER V0 ;
      RECT 1024 587 1056 619 ;
    LAYER V0 ;
      RECT 1024 587 1056 619 ;
    LAYER V0 ;
      RECT 1024 671 1056 703 ;
    LAYER V0 ;
      RECT 1024 671 1056 703 ;
    LAYER V0 ;
      RECT 1104 335 1136 367 ;
    LAYER V0 ;
      RECT 1104 419 1136 451 ;
    LAYER V0 ;
      RECT 1104 503 1136 535 ;
    LAYER V0 ;
      RECT 1104 587 1136 619 ;
    LAYER V0 ;
      RECT 1104 671 1136 703 ;
    LAYER V0 ;
      RECT 1104 908 1136 940 ;
    LAYER V0 ;
      RECT 1104 1748 1136 1780 ;
    LAYER V0 ;
      RECT 1184 335 1216 367 ;
    LAYER V0 ;
      RECT 1184 419 1216 451 ;
    LAYER V0 ;
      RECT 1184 503 1216 535 ;
    LAYER V0 ;
      RECT 1184 587 1216 619 ;
    LAYER V0 ;
      RECT 1184 671 1216 703 ;
  END
END DP_NMOS_B_40344802_X3_Y1
MACRO DP_NMOS_B_40344802_X1_Y3
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_40344802_X1_Y3 0 0 ;
  SIZE 800 BY 4704 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 4100 516 4132 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 60 48 100 2472 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 140 132 180 2556 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 220 888 260 3312 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 300 972 340 3396 ;
    END
  END GB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 380 216 420 2640 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1224 336 1968 ;
    LAYER M1 ;
      RECT 304 2064 336 2304 ;
    LAYER M1 ;
      RECT 304 2400 336 3144 ;
    LAYER M1 ;
      RECT 304 3240 336 3480 ;
    LAYER M1 ;
      RECT 304 3996 336 4236 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 224 1224 256 1968 ;
    LAYER M1 ;
      RECT 224 2400 256 3144 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 384 1224 416 1968 ;
    LAYER M1 ;
      RECT 384 2400 416 3144 ;
    LAYER M1 ;
      RECT 464 48 496 792 ;
    LAYER M1 ;
      RECT 464 888 496 1128 ;
    LAYER M1 ;
      RECT 464 1224 496 1968 ;
    LAYER M1 ;
      RECT 464 2064 496 2304 ;
    LAYER M1 ;
      RECT 464 2400 496 3144 ;
    LAYER M1 ;
      RECT 464 3240 496 3480 ;
    LAYER M1 ;
      RECT 464 3996 496 4236 ;
    LAYER M1 ;
      RECT 544 48 576 792 ;
    LAYER M1 ;
      RECT 544 1224 576 1968 ;
    LAYER M1 ;
      RECT 544 2400 576 3144 ;
    LAYER M2 ;
      RECT 44 68 356 100 ;
    LAYER M2 ;
      RECT 124 152 516 184 ;
    LAYER M2 ;
      RECT 124 908 356 940 ;
    LAYER M2 ;
      RECT 284 992 516 1024 ;
    LAYER M2 ;
      RECT 204 236 596 268 ;
    LAYER M2 ;
      RECT 44 1244 516 1276 ;
    LAYER M2 ;
      RECT 124 1328 356 1360 ;
    LAYER M2 ;
      RECT 204 2084 516 2116 ;
    LAYER M2 ;
      RECT 124 2168 356 2200 ;
    LAYER M2 ;
      RECT 204 1412 596 1444 ;
    LAYER M2 ;
      RECT 44 2420 356 2452 ;
    LAYER M2 ;
      RECT 124 2504 516 2536 ;
    LAYER M2 ;
      RECT 124 3260 356 3292 ;
    LAYER M2 ;
      RECT 284 3344 516 3376 ;
    LAYER M2 ;
      RECT 204 2588 596 2620 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1328 336 1360 ;
    LAYER V1 ;
      RECT 304 2168 336 2200 ;
    LAYER V1 ;
      RECT 304 2420 336 2452 ;
    LAYER V1 ;
      RECT 304 3260 336 3292 ;
    LAYER V1 ;
      RECT 304 4100 336 4132 ;
    LAYER V1 ;
      RECT 464 152 496 184 ;
    LAYER V1 ;
      RECT 464 992 496 1024 ;
    LAYER V1 ;
      RECT 464 1244 496 1276 ;
    LAYER V1 ;
      RECT 464 2084 496 2116 ;
    LAYER V1 ;
      RECT 464 2504 496 2536 ;
    LAYER V1 ;
      RECT 464 3344 496 3376 ;
    LAYER V1 ;
      RECT 464 4100 496 4132 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 224 1412 256 1444 ;
    LAYER V1 ;
      RECT 224 2588 256 2620 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 384 1412 416 1444 ;
    LAYER V1 ;
      RECT 384 2588 416 2620 ;
    LAYER V1 ;
      RECT 544 236 576 268 ;
    LAYER V1 ;
      RECT 544 1412 576 1444 ;
    LAYER V1 ;
      RECT 544 2588 576 2620 ;
    LAYER V2 ;
      RECT 64 68 96 100 ;
    LAYER V2 ;
      RECT 64 1244 96 1276 ;
    LAYER V2 ;
      RECT 64 2420 96 2452 ;
    LAYER V2 ;
      RECT 144 152 176 184 ;
    LAYER V2 ;
      RECT 144 1328 176 1360 ;
    LAYER V2 ;
      RECT 144 2504 176 2536 ;
    LAYER V2 ;
      RECT 224 908 256 940 ;
    LAYER V2 ;
      RECT 224 2084 256 2116 ;
    LAYER V2 ;
      RECT 224 3260 256 3292 ;
    LAYER V2 ;
      RECT 304 992 336 1024 ;
    LAYER V2 ;
      RECT 304 2168 336 2200 ;
    LAYER V2 ;
      RECT 304 3344 336 3376 ;
    LAYER V2 ;
      RECT 384 236 416 268 ;
    LAYER V2 ;
      RECT 384 1412 416 1444 ;
    LAYER V2 ;
      RECT 384 2588 416 2620 ;
    LAYER V0 ;
      RECT 304 335 336 367 ;
    LAYER V0 ;
      RECT 304 419 336 451 ;
    LAYER V0 ;
      RECT 304 503 336 535 ;
    LAYER V0 ;
      RECT 304 587 336 619 ;
    LAYER V0 ;
      RECT 304 671 336 703 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1511 336 1543 ;
    LAYER V0 ;
      RECT 304 1595 336 1627 ;
    LAYER V0 ;
      RECT 304 1679 336 1711 ;
    LAYER V0 ;
      RECT 304 1763 336 1795 ;
    LAYER V0 ;
      RECT 304 1847 336 1879 ;
    LAYER V0 ;
      RECT 304 2084 336 2116 ;
    LAYER V0 ;
      RECT 304 2687 336 2719 ;
    LAYER V0 ;
      RECT 304 2771 336 2803 ;
    LAYER V0 ;
      RECT 304 2855 336 2887 ;
    LAYER V0 ;
      RECT 304 2939 336 2971 ;
    LAYER V0 ;
      RECT 304 3023 336 3055 ;
    LAYER V0 ;
      RECT 304 3260 336 3292 ;
    LAYER V0 ;
      RECT 304 4100 336 4132 ;
    LAYER V0 ;
      RECT 304 4100 336 4132 ;
    LAYER V0 ;
      RECT 304 4100 336 4132 ;
    LAYER V0 ;
      RECT 224 335 256 367 ;
    LAYER V0 ;
      RECT 224 419 256 451 ;
    LAYER V0 ;
      RECT 224 503 256 535 ;
    LAYER V0 ;
      RECT 224 587 256 619 ;
    LAYER V0 ;
      RECT 224 671 256 703 ;
    LAYER V0 ;
      RECT 224 1511 256 1543 ;
    LAYER V0 ;
      RECT 224 1595 256 1627 ;
    LAYER V0 ;
      RECT 224 1679 256 1711 ;
    LAYER V0 ;
      RECT 224 1763 256 1795 ;
    LAYER V0 ;
      RECT 224 1847 256 1879 ;
    LAYER V0 ;
      RECT 224 2687 256 2719 ;
    LAYER V0 ;
      RECT 224 2771 256 2803 ;
    LAYER V0 ;
      RECT 224 2855 256 2887 ;
    LAYER V0 ;
      RECT 224 2939 256 2971 ;
    LAYER V0 ;
      RECT 224 3023 256 3055 ;
    LAYER V0 ;
      RECT 384 335 416 367 ;
    LAYER V0 ;
      RECT 384 335 416 367 ;
    LAYER V0 ;
      RECT 384 419 416 451 ;
    LAYER V0 ;
      RECT 384 419 416 451 ;
    LAYER V0 ;
      RECT 384 503 416 535 ;
    LAYER V0 ;
      RECT 384 503 416 535 ;
    LAYER V0 ;
      RECT 384 587 416 619 ;
    LAYER V0 ;
      RECT 384 587 416 619 ;
    LAYER V0 ;
      RECT 384 671 416 703 ;
    LAYER V0 ;
      RECT 384 671 416 703 ;
    LAYER V0 ;
      RECT 384 1511 416 1543 ;
    LAYER V0 ;
      RECT 384 1511 416 1543 ;
    LAYER V0 ;
      RECT 384 1595 416 1627 ;
    LAYER V0 ;
      RECT 384 1595 416 1627 ;
    LAYER V0 ;
      RECT 384 1679 416 1711 ;
    LAYER V0 ;
      RECT 384 1679 416 1711 ;
    LAYER V0 ;
      RECT 384 1763 416 1795 ;
    LAYER V0 ;
      RECT 384 1763 416 1795 ;
    LAYER V0 ;
      RECT 384 1847 416 1879 ;
    LAYER V0 ;
      RECT 384 1847 416 1879 ;
    LAYER V0 ;
      RECT 384 2687 416 2719 ;
    LAYER V0 ;
      RECT 384 2687 416 2719 ;
    LAYER V0 ;
      RECT 384 2771 416 2803 ;
    LAYER V0 ;
      RECT 384 2771 416 2803 ;
    LAYER V0 ;
      RECT 384 2855 416 2887 ;
    LAYER V0 ;
      RECT 384 2855 416 2887 ;
    LAYER V0 ;
      RECT 384 2939 416 2971 ;
    LAYER V0 ;
      RECT 384 2939 416 2971 ;
    LAYER V0 ;
      RECT 384 3023 416 3055 ;
    LAYER V0 ;
      RECT 384 3023 416 3055 ;
    LAYER V0 ;
      RECT 464 335 496 367 ;
    LAYER V0 ;
      RECT 464 419 496 451 ;
    LAYER V0 ;
      RECT 464 503 496 535 ;
    LAYER V0 ;
      RECT 464 587 496 619 ;
    LAYER V0 ;
      RECT 464 671 496 703 ;
    LAYER V0 ;
      RECT 464 908 496 940 ;
    LAYER V0 ;
      RECT 464 1511 496 1543 ;
    LAYER V0 ;
      RECT 464 1595 496 1627 ;
    LAYER V0 ;
      RECT 464 1679 496 1711 ;
    LAYER V0 ;
      RECT 464 1763 496 1795 ;
    LAYER V0 ;
      RECT 464 1847 496 1879 ;
    LAYER V0 ;
      RECT 464 2084 496 2116 ;
    LAYER V0 ;
      RECT 464 2687 496 2719 ;
    LAYER V0 ;
      RECT 464 2771 496 2803 ;
    LAYER V0 ;
      RECT 464 2855 496 2887 ;
    LAYER V0 ;
      RECT 464 2939 496 2971 ;
    LAYER V0 ;
      RECT 464 3023 496 3055 ;
    LAYER V0 ;
      RECT 464 3260 496 3292 ;
    LAYER V0 ;
      RECT 464 4100 496 4132 ;
    LAYER V0 ;
      RECT 464 4100 496 4132 ;
    LAYER V0 ;
      RECT 464 4100 496 4132 ;
    LAYER V0 ;
      RECT 544 335 576 367 ;
    LAYER V0 ;
      RECT 544 419 576 451 ;
    LAYER V0 ;
      RECT 544 503 576 535 ;
    LAYER V0 ;
      RECT 544 587 576 619 ;
    LAYER V0 ;
      RECT 544 671 576 703 ;
    LAYER V0 ;
      RECT 544 1511 576 1543 ;
    LAYER V0 ;
      RECT 544 1595 576 1627 ;
    LAYER V0 ;
      RECT 544 1679 576 1711 ;
    LAYER V0 ;
      RECT 544 1763 576 1795 ;
    LAYER V0 ;
      RECT 544 1847 576 1879 ;
    LAYER V0 ;
      RECT 544 2687 576 2719 ;
    LAYER V0 ;
      RECT 544 2771 576 2803 ;
    LAYER V0 ;
      RECT 544 2855 576 2887 ;
    LAYER V0 ;
      RECT 544 2939 576 2971 ;
    LAYER V0 ;
      RECT 544 3023 576 3055 ;
  END
END DP_NMOS_B_40344802_X1_Y3
MACRO CAP_12F
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CAP_12F 0 0 ;
  SIZE 8400 BY 8148 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44 7964 8356 7996 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44 152 8356 184 ;
    END
  END PLUS
  OBS
    LAYER M1 ;
      RECT 304 132 336 8016 ;
    LAYER M1 ;
      RECT 368 132 400 8016 ;
    LAYER M1 ;
      RECT 432 132 464 8016 ;
    LAYER M1 ;
      RECT 496 132 528 8016 ;
    LAYER M1 ;
      RECT 560 132 592 8016 ;
    LAYER M1 ;
      RECT 624 132 656 8016 ;
    LAYER M1 ;
      RECT 688 132 720 8016 ;
    LAYER M1 ;
      RECT 752 132 784 8016 ;
    LAYER M1 ;
      RECT 816 132 848 8016 ;
    LAYER M1 ;
      RECT 880 132 912 8016 ;
    LAYER M1 ;
      RECT 944 132 976 8016 ;
    LAYER M1 ;
      RECT 1008 132 1040 8016 ;
    LAYER M1 ;
      RECT 1072 132 1104 8016 ;
    LAYER M1 ;
      RECT 1136 132 1168 8016 ;
    LAYER M1 ;
      RECT 1200 132 1232 8016 ;
    LAYER M1 ;
      RECT 1264 132 1296 8016 ;
    LAYER M1 ;
      RECT 1328 132 1360 8016 ;
    LAYER M1 ;
      RECT 1392 132 1424 8016 ;
    LAYER M1 ;
      RECT 1456 132 1488 8016 ;
    LAYER M1 ;
      RECT 1520 132 1552 8016 ;
    LAYER M1 ;
      RECT 1584 132 1616 8016 ;
    LAYER M1 ;
      RECT 1648 132 1680 8016 ;
    LAYER M1 ;
      RECT 1712 132 1744 8016 ;
    LAYER M1 ;
      RECT 1776 132 1808 8016 ;
    LAYER M1 ;
      RECT 1840 132 1872 8016 ;
    LAYER M1 ;
      RECT 1904 132 1936 8016 ;
    LAYER M1 ;
      RECT 1968 132 2000 8016 ;
    LAYER M1 ;
      RECT 2032 132 2064 8016 ;
    LAYER M1 ;
      RECT 2096 132 2128 8016 ;
    LAYER M1 ;
      RECT 2160 132 2192 8016 ;
    LAYER M1 ;
      RECT 2224 132 2256 8016 ;
    LAYER M1 ;
      RECT 2288 132 2320 8016 ;
    LAYER M1 ;
      RECT 2352 132 2384 8016 ;
    LAYER M1 ;
      RECT 2416 132 2448 8016 ;
    LAYER M1 ;
      RECT 2480 132 2512 8016 ;
    LAYER M1 ;
      RECT 2544 132 2576 8016 ;
    LAYER M1 ;
      RECT 2608 132 2640 8016 ;
    LAYER M1 ;
      RECT 2672 132 2704 8016 ;
    LAYER M1 ;
      RECT 2736 132 2768 8016 ;
    LAYER M1 ;
      RECT 2800 132 2832 8016 ;
    LAYER M1 ;
      RECT 2864 132 2896 8016 ;
    LAYER M1 ;
      RECT 2928 132 2960 8016 ;
    LAYER M1 ;
      RECT 2992 132 3024 8016 ;
    LAYER M1 ;
      RECT 3056 132 3088 8016 ;
    LAYER M1 ;
      RECT 3120 132 3152 8016 ;
    LAYER M1 ;
      RECT 3184 132 3216 8016 ;
    LAYER M1 ;
      RECT 3248 132 3280 8016 ;
    LAYER M1 ;
      RECT 3312 132 3344 8016 ;
    LAYER M1 ;
      RECT 3376 132 3408 8016 ;
    LAYER M1 ;
      RECT 3440 132 3472 8016 ;
    LAYER M1 ;
      RECT 3504 132 3536 8016 ;
    LAYER M1 ;
      RECT 3568 132 3600 8016 ;
    LAYER M1 ;
      RECT 3632 132 3664 8016 ;
    LAYER M1 ;
      RECT 3696 132 3728 8016 ;
    LAYER M1 ;
      RECT 3760 132 3792 8016 ;
    LAYER M1 ;
      RECT 3824 132 3856 8016 ;
    LAYER M1 ;
      RECT 3888 132 3920 8016 ;
    LAYER M1 ;
      RECT 3952 132 3984 8016 ;
    LAYER M1 ;
      RECT 4016 132 4048 8016 ;
    LAYER M1 ;
      RECT 4080 132 4112 8016 ;
    LAYER M1 ;
      RECT 4144 132 4176 8016 ;
    LAYER M1 ;
      RECT 4208 132 4240 8016 ;
    LAYER M1 ;
      RECT 4272 132 4304 8016 ;
    LAYER M1 ;
      RECT 4336 132 4368 8016 ;
    LAYER M1 ;
      RECT 4400 132 4432 8016 ;
    LAYER M1 ;
      RECT 4464 132 4496 8016 ;
    LAYER M1 ;
      RECT 4528 132 4560 8016 ;
    LAYER M1 ;
      RECT 4592 132 4624 8016 ;
    LAYER M1 ;
      RECT 4656 132 4688 8016 ;
    LAYER M1 ;
      RECT 4720 132 4752 8016 ;
    LAYER M1 ;
      RECT 4784 132 4816 8016 ;
    LAYER M1 ;
      RECT 4848 132 4880 8016 ;
    LAYER M1 ;
      RECT 4912 132 4944 8016 ;
    LAYER M1 ;
      RECT 4976 132 5008 8016 ;
    LAYER M1 ;
      RECT 5040 132 5072 8016 ;
    LAYER M1 ;
      RECT 5104 132 5136 8016 ;
    LAYER M1 ;
      RECT 5168 132 5200 8016 ;
    LAYER M1 ;
      RECT 5232 132 5264 8016 ;
    LAYER M1 ;
      RECT 5296 132 5328 8016 ;
    LAYER M1 ;
      RECT 5360 132 5392 8016 ;
    LAYER M1 ;
      RECT 5424 132 5456 8016 ;
    LAYER M1 ;
      RECT 5488 132 5520 8016 ;
    LAYER M1 ;
      RECT 5552 132 5584 8016 ;
    LAYER M1 ;
      RECT 5616 132 5648 8016 ;
    LAYER M1 ;
      RECT 5680 132 5712 8016 ;
    LAYER M1 ;
      RECT 5744 132 5776 8016 ;
    LAYER M1 ;
      RECT 5808 132 5840 8016 ;
    LAYER M1 ;
      RECT 5872 132 5904 8016 ;
    LAYER M1 ;
      RECT 5936 132 5968 8016 ;
    LAYER M1 ;
      RECT 6000 132 6032 8016 ;
    LAYER M1 ;
      RECT 6064 132 6096 8016 ;
    LAYER M1 ;
      RECT 6128 132 6160 8016 ;
    LAYER M1 ;
      RECT 6192 132 6224 8016 ;
    LAYER M1 ;
      RECT 6256 132 6288 8016 ;
    LAYER M1 ;
      RECT 6320 132 6352 8016 ;
    LAYER M1 ;
      RECT 6384 132 6416 8016 ;
    LAYER M1 ;
      RECT 6448 132 6480 8016 ;
    LAYER M1 ;
      RECT 6512 132 6544 8016 ;
    LAYER M1 ;
      RECT 6576 132 6608 8016 ;
    LAYER M1 ;
      RECT 6640 132 6672 8016 ;
    LAYER M1 ;
      RECT 6704 132 6736 8016 ;
    LAYER M1 ;
      RECT 6768 132 6800 8016 ;
    LAYER M1 ;
      RECT 6832 132 6864 8016 ;
    LAYER M1 ;
      RECT 6896 132 6928 8016 ;
    LAYER M1 ;
      RECT 6960 132 6992 8016 ;
    LAYER M1 ;
      RECT 7024 132 7056 8016 ;
    LAYER M1 ;
      RECT 7088 132 7120 8016 ;
    LAYER M1 ;
      RECT 7152 132 7184 8016 ;
    LAYER M1 ;
      RECT 7216 132 7248 8016 ;
    LAYER M1 ;
      RECT 7280 132 7312 8016 ;
    LAYER M1 ;
      RECT 7344 132 7376 8016 ;
    LAYER M1 ;
      RECT 7408 132 7440 8016 ;
    LAYER M1 ;
      RECT 7472 132 7504 8016 ;
    LAYER M1 ;
      RECT 7536 132 7568 8016 ;
    LAYER M1 ;
      RECT 7600 132 7632 8016 ;
    LAYER M1 ;
      RECT 7664 132 7696 8016 ;
    LAYER M1 ;
      RECT 7728 132 7760 8016 ;
    LAYER M1 ;
      RECT 7792 132 7824 8016 ;
    LAYER M1 ;
      RECT 7856 132 7888 8016 ;
    LAYER M1 ;
      RECT 7920 132 7952 8016 ;
    LAYER M1 ;
      RECT 7984 132 8016 8016 ;
    LAYER M1 ;
      RECT 8064 132 8096 8016 ;
    LAYER M2 ;
      RECT 284 216 8116 248 ;
    LAYER M2 ;
      RECT 284 280 8116 312 ;
    LAYER M2 ;
      RECT 284 344 8116 376 ;
    LAYER M2 ;
      RECT 284 408 8116 440 ;
    LAYER M2 ;
      RECT 284 472 8116 504 ;
    LAYER M2 ;
      RECT 284 536 8116 568 ;
    LAYER M2 ;
      RECT 284 600 8116 632 ;
    LAYER M2 ;
      RECT 284 664 8116 696 ;
    LAYER M2 ;
      RECT 284 728 8116 760 ;
    LAYER M2 ;
      RECT 284 792 8116 824 ;
    LAYER M2 ;
      RECT 284 856 8116 888 ;
    LAYER M2 ;
      RECT 284 920 8116 952 ;
    LAYER M2 ;
      RECT 284 984 8116 1016 ;
    LAYER M2 ;
      RECT 284 1048 8116 1080 ;
    LAYER M2 ;
      RECT 284 1112 8116 1144 ;
    LAYER M2 ;
      RECT 284 1176 8116 1208 ;
    LAYER M2 ;
      RECT 284 1240 8116 1272 ;
    LAYER M2 ;
      RECT 284 1304 8116 1336 ;
    LAYER M2 ;
      RECT 284 1368 8116 1400 ;
    LAYER M2 ;
      RECT 284 1432 8116 1464 ;
    LAYER M2 ;
      RECT 284 1496 8116 1528 ;
    LAYER M2 ;
      RECT 284 1560 8116 1592 ;
    LAYER M2 ;
      RECT 284 1624 8116 1656 ;
    LAYER M2 ;
      RECT 284 1688 8116 1720 ;
    LAYER M2 ;
      RECT 284 1752 8116 1784 ;
    LAYER M2 ;
      RECT 284 1816 8116 1848 ;
    LAYER M2 ;
      RECT 284 1880 8116 1912 ;
    LAYER M2 ;
      RECT 284 1944 8116 1976 ;
    LAYER M2 ;
      RECT 284 2008 8116 2040 ;
    LAYER M2 ;
      RECT 284 2072 8116 2104 ;
    LAYER M2 ;
      RECT 284 2136 8116 2168 ;
    LAYER M2 ;
      RECT 284 2200 8116 2232 ;
    LAYER M2 ;
      RECT 284 2264 8116 2296 ;
    LAYER M2 ;
      RECT 284 2328 8116 2360 ;
    LAYER M2 ;
      RECT 284 2392 8116 2424 ;
    LAYER M2 ;
      RECT 284 2456 8116 2488 ;
    LAYER M2 ;
      RECT 284 2520 8116 2552 ;
    LAYER M2 ;
      RECT 284 2584 8116 2616 ;
    LAYER M2 ;
      RECT 284 2648 8116 2680 ;
    LAYER M2 ;
      RECT 284 2712 8116 2744 ;
    LAYER M2 ;
      RECT 284 2776 8116 2808 ;
    LAYER M2 ;
      RECT 284 2840 8116 2872 ;
    LAYER M2 ;
      RECT 284 2904 8116 2936 ;
    LAYER M2 ;
      RECT 284 2968 8116 3000 ;
    LAYER M2 ;
      RECT 284 3032 8116 3064 ;
    LAYER M2 ;
      RECT 284 3096 8116 3128 ;
    LAYER M2 ;
      RECT 284 3160 8116 3192 ;
    LAYER M2 ;
      RECT 284 3224 8116 3256 ;
    LAYER M2 ;
      RECT 284 3288 8116 3320 ;
    LAYER M2 ;
      RECT 284 3352 8116 3384 ;
    LAYER M2 ;
      RECT 284 3416 8116 3448 ;
    LAYER M2 ;
      RECT 284 3480 8116 3512 ;
    LAYER M2 ;
      RECT 284 3544 8116 3576 ;
    LAYER M2 ;
      RECT 284 3608 8116 3640 ;
    LAYER M2 ;
      RECT 284 3672 8116 3704 ;
    LAYER M2 ;
      RECT 284 3736 8116 3768 ;
    LAYER M2 ;
      RECT 284 3800 8116 3832 ;
    LAYER M2 ;
      RECT 284 3864 8116 3896 ;
    LAYER M2 ;
      RECT 284 3928 8116 3960 ;
    LAYER M2 ;
      RECT 284 3992 8116 4024 ;
    LAYER M2 ;
      RECT 284 4056 8116 4088 ;
    LAYER M2 ;
      RECT 284 4120 8116 4152 ;
    LAYER M2 ;
      RECT 284 4184 8116 4216 ;
    LAYER M2 ;
      RECT 284 4248 8116 4280 ;
    LAYER M2 ;
      RECT 284 4312 8116 4344 ;
    LAYER M2 ;
      RECT 284 4376 8116 4408 ;
    LAYER M2 ;
      RECT 284 4440 8116 4472 ;
    LAYER M2 ;
      RECT 284 4504 8116 4536 ;
    LAYER M2 ;
      RECT 284 4568 8116 4600 ;
    LAYER M2 ;
      RECT 284 4632 8116 4664 ;
    LAYER M2 ;
      RECT 284 4696 8116 4728 ;
    LAYER M2 ;
      RECT 284 4760 8116 4792 ;
    LAYER M2 ;
      RECT 284 4824 8116 4856 ;
    LAYER M2 ;
      RECT 284 4888 8116 4920 ;
    LAYER M2 ;
      RECT 284 4952 8116 4984 ;
    LAYER M2 ;
      RECT 284 5016 8116 5048 ;
    LAYER M2 ;
      RECT 284 5080 8116 5112 ;
    LAYER M2 ;
      RECT 284 5144 8116 5176 ;
    LAYER M2 ;
      RECT 284 5208 8116 5240 ;
    LAYER M2 ;
      RECT 284 5272 8116 5304 ;
    LAYER M2 ;
      RECT 284 5336 8116 5368 ;
    LAYER M2 ;
      RECT 284 5400 8116 5432 ;
    LAYER M2 ;
      RECT 284 5464 8116 5496 ;
    LAYER M2 ;
      RECT 284 5528 8116 5560 ;
    LAYER M2 ;
      RECT 284 5592 8116 5624 ;
    LAYER M2 ;
      RECT 284 5656 8116 5688 ;
    LAYER M2 ;
      RECT 284 5720 8116 5752 ;
    LAYER M2 ;
      RECT 284 5784 8116 5816 ;
    LAYER M2 ;
      RECT 284 5848 8116 5880 ;
    LAYER M2 ;
      RECT 284 5912 8116 5944 ;
    LAYER M2 ;
      RECT 284 5976 8116 6008 ;
    LAYER M2 ;
      RECT 284 6040 8116 6072 ;
    LAYER M2 ;
      RECT 284 6104 8116 6136 ;
    LAYER M2 ;
      RECT 284 6168 8116 6200 ;
    LAYER M2 ;
      RECT 284 6232 8116 6264 ;
    LAYER M2 ;
      RECT 284 6296 8116 6328 ;
    LAYER M2 ;
      RECT 284 6360 8116 6392 ;
    LAYER M2 ;
      RECT 284 6424 8116 6456 ;
    LAYER M2 ;
      RECT 284 6488 8116 6520 ;
    LAYER M2 ;
      RECT 284 6552 8116 6584 ;
    LAYER M2 ;
      RECT 284 6616 8116 6648 ;
    LAYER M2 ;
      RECT 284 6680 8116 6712 ;
    LAYER M2 ;
      RECT 284 6744 8116 6776 ;
    LAYER M2 ;
      RECT 284 6808 8116 6840 ;
    LAYER M2 ;
      RECT 284 6872 8116 6904 ;
    LAYER M2 ;
      RECT 284 6936 8116 6968 ;
    LAYER M2 ;
      RECT 284 7000 8116 7032 ;
    LAYER M2 ;
      RECT 284 7064 8116 7096 ;
    LAYER M2 ;
      RECT 284 7128 8116 7160 ;
    LAYER M2 ;
      RECT 284 7192 8116 7224 ;
    LAYER M2 ;
      RECT 284 7256 8116 7288 ;
    LAYER M2 ;
      RECT 284 7320 8116 7352 ;
    LAYER M2 ;
      RECT 284 7384 8116 7416 ;
    LAYER M2 ;
      RECT 284 7448 8116 7480 ;
    LAYER M2 ;
      RECT 284 7512 8116 7544 ;
    LAYER M2 ;
      RECT 284 7576 8116 7608 ;
    LAYER M2 ;
      RECT 284 7640 8116 7672 ;
    LAYER M2 ;
      RECT 284 7704 8116 7736 ;
    LAYER M2 ;
      RECT 284 7768 8116 7800 ;
    LAYER M2 ;
      RECT 284 7832 8116 7864 ;
    LAYER V1 ;
      RECT 304 216 336 248 ;
    LAYER V1 ;
      RECT 304 344 336 376 ;
    LAYER V1 ;
      RECT 304 472 336 504 ;
    LAYER V1 ;
      RECT 304 600 336 632 ;
    LAYER V1 ;
      RECT 304 728 336 760 ;
    LAYER V1 ;
      RECT 304 856 336 888 ;
    LAYER V1 ;
      RECT 304 984 336 1016 ;
    LAYER V1 ;
      RECT 304 1112 336 1144 ;
    LAYER V1 ;
      RECT 304 1240 336 1272 ;
    LAYER V1 ;
      RECT 304 1368 336 1400 ;
    LAYER V1 ;
      RECT 304 1496 336 1528 ;
    LAYER V1 ;
      RECT 304 1624 336 1656 ;
    LAYER V1 ;
      RECT 304 1752 336 1784 ;
    LAYER V1 ;
      RECT 304 1880 336 1912 ;
    LAYER V1 ;
      RECT 304 2008 336 2040 ;
    LAYER V1 ;
      RECT 304 2136 336 2168 ;
    LAYER V1 ;
      RECT 304 2264 336 2296 ;
    LAYER V1 ;
      RECT 304 2392 336 2424 ;
    LAYER V1 ;
      RECT 304 2520 336 2552 ;
    LAYER V1 ;
      RECT 304 2648 336 2680 ;
    LAYER V1 ;
      RECT 304 2776 336 2808 ;
    LAYER V1 ;
      RECT 304 2904 336 2936 ;
    LAYER V1 ;
      RECT 304 3032 336 3064 ;
    LAYER V1 ;
      RECT 304 3160 336 3192 ;
    LAYER V1 ;
      RECT 304 3288 336 3320 ;
    LAYER V1 ;
      RECT 304 3416 336 3448 ;
    LAYER V1 ;
      RECT 304 3544 336 3576 ;
    LAYER V1 ;
      RECT 304 3672 336 3704 ;
    LAYER V1 ;
      RECT 304 3800 336 3832 ;
    LAYER V1 ;
      RECT 304 3928 336 3960 ;
    LAYER V1 ;
      RECT 304 4056 336 4088 ;
    LAYER V1 ;
      RECT 304 4184 336 4216 ;
    LAYER V1 ;
      RECT 304 4312 336 4344 ;
    LAYER V1 ;
      RECT 304 4440 336 4472 ;
    LAYER V1 ;
      RECT 304 4568 336 4600 ;
    LAYER V1 ;
      RECT 304 4696 336 4728 ;
    LAYER V1 ;
      RECT 304 4824 336 4856 ;
    LAYER V1 ;
      RECT 304 4952 336 4984 ;
    LAYER V1 ;
      RECT 304 5080 336 5112 ;
    LAYER V1 ;
      RECT 304 5208 336 5240 ;
    LAYER V1 ;
      RECT 304 5336 336 5368 ;
    LAYER V1 ;
      RECT 304 5464 336 5496 ;
    LAYER V1 ;
      RECT 304 5592 336 5624 ;
    LAYER V1 ;
      RECT 304 5720 336 5752 ;
    LAYER V1 ;
      RECT 304 5848 336 5880 ;
    LAYER V1 ;
      RECT 304 5976 336 6008 ;
    LAYER V1 ;
      RECT 304 6104 336 6136 ;
    LAYER V1 ;
      RECT 304 6232 336 6264 ;
    LAYER V1 ;
      RECT 304 6360 336 6392 ;
    LAYER V1 ;
      RECT 304 6488 336 6520 ;
    LAYER V1 ;
      RECT 304 6616 336 6648 ;
    LAYER V1 ;
      RECT 304 6744 336 6776 ;
    LAYER V1 ;
      RECT 304 6872 336 6904 ;
    LAYER V1 ;
      RECT 304 7000 336 7032 ;
    LAYER V1 ;
      RECT 304 7128 336 7160 ;
    LAYER V1 ;
      RECT 304 7256 336 7288 ;
    LAYER V1 ;
      RECT 304 7384 336 7416 ;
    LAYER V1 ;
      RECT 304 7512 336 7544 ;
    LAYER V1 ;
      RECT 304 7640 336 7672 ;
    LAYER V1 ;
      RECT 304 7768 336 7800 ;
    LAYER V1 ;
      RECT 304 7964 336 7996 ;
    LAYER V1 ;
      RECT 368 152 400 184 ;
    LAYER V1 ;
      RECT 432 7964 464 7996 ;
    LAYER V1 ;
      RECT 496 152 528 184 ;
    LAYER V1 ;
      RECT 560 7964 592 7996 ;
    LAYER V1 ;
      RECT 624 152 656 184 ;
    LAYER V1 ;
      RECT 688 7964 720 7996 ;
    LAYER V1 ;
      RECT 752 152 784 184 ;
    LAYER V1 ;
      RECT 816 7964 848 7996 ;
    LAYER V1 ;
      RECT 880 152 912 184 ;
    LAYER V1 ;
      RECT 944 7964 976 7996 ;
    LAYER V1 ;
      RECT 1008 152 1040 184 ;
    LAYER V1 ;
      RECT 1072 7964 1104 7996 ;
    LAYER V1 ;
      RECT 1136 152 1168 184 ;
    LAYER V1 ;
      RECT 1200 7964 1232 7996 ;
    LAYER V1 ;
      RECT 1264 152 1296 184 ;
    LAYER V1 ;
      RECT 1328 7964 1360 7996 ;
    LAYER V1 ;
      RECT 1392 152 1424 184 ;
    LAYER V1 ;
      RECT 1456 7964 1488 7996 ;
    LAYER V1 ;
      RECT 1520 152 1552 184 ;
    LAYER V1 ;
      RECT 1584 7964 1616 7996 ;
    LAYER V1 ;
      RECT 1648 152 1680 184 ;
    LAYER V1 ;
      RECT 1712 7964 1744 7996 ;
    LAYER V1 ;
      RECT 1776 152 1808 184 ;
    LAYER V1 ;
      RECT 1840 7964 1872 7996 ;
    LAYER V1 ;
      RECT 1904 152 1936 184 ;
    LAYER V1 ;
      RECT 1968 7964 2000 7996 ;
    LAYER V1 ;
      RECT 2032 152 2064 184 ;
    LAYER V1 ;
      RECT 2096 7964 2128 7996 ;
    LAYER V1 ;
      RECT 2160 152 2192 184 ;
    LAYER V1 ;
      RECT 2224 7964 2256 7996 ;
    LAYER V1 ;
      RECT 2288 152 2320 184 ;
    LAYER V1 ;
      RECT 2352 7964 2384 7996 ;
    LAYER V1 ;
      RECT 2416 152 2448 184 ;
    LAYER V1 ;
      RECT 2480 7964 2512 7996 ;
    LAYER V1 ;
      RECT 2544 152 2576 184 ;
    LAYER V1 ;
      RECT 2608 7964 2640 7996 ;
    LAYER V1 ;
      RECT 2672 152 2704 184 ;
    LAYER V1 ;
      RECT 2736 7964 2768 7996 ;
    LAYER V1 ;
      RECT 2800 152 2832 184 ;
    LAYER V1 ;
      RECT 2864 7964 2896 7996 ;
    LAYER V1 ;
      RECT 2928 152 2960 184 ;
    LAYER V1 ;
      RECT 2992 7964 3024 7996 ;
    LAYER V1 ;
      RECT 3056 152 3088 184 ;
    LAYER V1 ;
      RECT 3120 7964 3152 7996 ;
    LAYER V1 ;
      RECT 3184 152 3216 184 ;
    LAYER V1 ;
      RECT 3248 7964 3280 7996 ;
    LAYER V1 ;
      RECT 3312 152 3344 184 ;
    LAYER V1 ;
      RECT 3376 7964 3408 7996 ;
    LAYER V1 ;
      RECT 3440 152 3472 184 ;
    LAYER V1 ;
      RECT 3504 7964 3536 7996 ;
    LAYER V1 ;
      RECT 3568 152 3600 184 ;
    LAYER V1 ;
      RECT 3632 7964 3664 7996 ;
    LAYER V1 ;
      RECT 3696 152 3728 184 ;
    LAYER V1 ;
      RECT 3760 7964 3792 7996 ;
    LAYER V1 ;
      RECT 3824 152 3856 184 ;
    LAYER V1 ;
      RECT 3888 7964 3920 7996 ;
    LAYER V1 ;
      RECT 3952 152 3984 184 ;
    LAYER V1 ;
      RECT 4016 7964 4048 7996 ;
    LAYER V1 ;
      RECT 4080 152 4112 184 ;
    LAYER V1 ;
      RECT 4144 7964 4176 7996 ;
    LAYER V1 ;
      RECT 4208 152 4240 184 ;
    LAYER V1 ;
      RECT 4272 7964 4304 7996 ;
    LAYER V1 ;
      RECT 4336 152 4368 184 ;
    LAYER V1 ;
      RECT 4400 7964 4432 7996 ;
    LAYER V1 ;
      RECT 4464 152 4496 184 ;
    LAYER V1 ;
      RECT 4528 7964 4560 7996 ;
    LAYER V1 ;
      RECT 4592 152 4624 184 ;
    LAYER V1 ;
      RECT 4656 7964 4688 7996 ;
    LAYER V1 ;
      RECT 4720 152 4752 184 ;
    LAYER V1 ;
      RECT 4784 7964 4816 7996 ;
    LAYER V1 ;
      RECT 4848 152 4880 184 ;
    LAYER V1 ;
      RECT 4912 7964 4944 7996 ;
    LAYER V1 ;
      RECT 4976 152 5008 184 ;
    LAYER V1 ;
      RECT 5040 7964 5072 7996 ;
    LAYER V1 ;
      RECT 5104 152 5136 184 ;
    LAYER V1 ;
      RECT 5168 7964 5200 7996 ;
    LAYER V1 ;
      RECT 5232 152 5264 184 ;
    LAYER V1 ;
      RECT 5296 7964 5328 7996 ;
    LAYER V1 ;
      RECT 5360 152 5392 184 ;
    LAYER V1 ;
      RECT 5424 7964 5456 7996 ;
    LAYER V1 ;
      RECT 5488 152 5520 184 ;
    LAYER V1 ;
      RECT 5552 7964 5584 7996 ;
    LAYER V1 ;
      RECT 5616 152 5648 184 ;
    LAYER V1 ;
      RECT 5680 7964 5712 7996 ;
    LAYER V1 ;
      RECT 5744 152 5776 184 ;
    LAYER V1 ;
      RECT 5808 7964 5840 7996 ;
    LAYER V1 ;
      RECT 5872 152 5904 184 ;
    LAYER V1 ;
      RECT 5936 7964 5968 7996 ;
    LAYER V1 ;
      RECT 6000 152 6032 184 ;
    LAYER V1 ;
      RECT 6064 7964 6096 7996 ;
    LAYER V1 ;
      RECT 6128 152 6160 184 ;
    LAYER V1 ;
      RECT 6192 7964 6224 7996 ;
    LAYER V1 ;
      RECT 6256 152 6288 184 ;
    LAYER V1 ;
      RECT 6320 7964 6352 7996 ;
    LAYER V1 ;
      RECT 6384 152 6416 184 ;
    LAYER V1 ;
      RECT 6448 7964 6480 7996 ;
    LAYER V1 ;
      RECT 6512 152 6544 184 ;
    LAYER V1 ;
      RECT 6576 7964 6608 7996 ;
    LAYER V1 ;
      RECT 6640 152 6672 184 ;
    LAYER V1 ;
      RECT 6704 7964 6736 7996 ;
    LAYER V1 ;
      RECT 6768 152 6800 184 ;
    LAYER V1 ;
      RECT 6832 7964 6864 7996 ;
    LAYER V1 ;
      RECT 6896 152 6928 184 ;
    LAYER V1 ;
      RECT 6960 7964 6992 7996 ;
    LAYER V1 ;
      RECT 7024 152 7056 184 ;
    LAYER V1 ;
      RECT 7088 7964 7120 7996 ;
    LAYER V1 ;
      RECT 7152 152 7184 184 ;
    LAYER V1 ;
      RECT 7216 7964 7248 7996 ;
    LAYER V1 ;
      RECT 7280 152 7312 184 ;
    LAYER V1 ;
      RECT 7344 7964 7376 7996 ;
    LAYER V1 ;
      RECT 7408 152 7440 184 ;
    LAYER V1 ;
      RECT 7472 7964 7504 7996 ;
    LAYER V1 ;
      RECT 7536 152 7568 184 ;
    LAYER V1 ;
      RECT 7600 7964 7632 7996 ;
    LAYER V1 ;
      RECT 7664 152 7696 184 ;
    LAYER V1 ;
      RECT 7728 7964 7760 7996 ;
    LAYER V1 ;
      RECT 7792 152 7824 184 ;
    LAYER V1 ;
      RECT 7856 7964 7888 7996 ;
    LAYER V1 ;
      RECT 7920 152 7952 184 ;
    LAYER V1 ;
      RECT 7984 7964 8016 7996 ;
    LAYER V1 ;
      RECT 8064 152 8096 184 ;
    LAYER V1 ;
      RECT 8064 280 8096 312 ;
    LAYER V1 ;
      RECT 8064 408 8096 440 ;
    LAYER V1 ;
      RECT 8064 536 8096 568 ;
    LAYER V1 ;
      RECT 8064 664 8096 696 ;
    LAYER V1 ;
      RECT 8064 792 8096 824 ;
    LAYER V1 ;
      RECT 8064 920 8096 952 ;
    LAYER V1 ;
      RECT 8064 1048 8096 1080 ;
    LAYER V1 ;
      RECT 8064 1176 8096 1208 ;
    LAYER V1 ;
      RECT 8064 1304 8096 1336 ;
    LAYER V1 ;
      RECT 8064 1432 8096 1464 ;
    LAYER V1 ;
      RECT 8064 1560 8096 1592 ;
    LAYER V1 ;
      RECT 8064 1688 8096 1720 ;
    LAYER V1 ;
      RECT 8064 1816 8096 1848 ;
    LAYER V1 ;
      RECT 8064 1944 8096 1976 ;
    LAYER V1 ;
      RECT 8064 2072 8096 2104 ;
    LAYER V1 ;
      RECT 8064 2200 8096 2232 ;
    LAYER V1 ;
      RECT 8064 2328 8096 2360 ;
    LAYER V1 ;
      RECT 8064 2456 8096 2488 ;
    LAYER V1 ;
      RECT 8064 2584 8096 2616 ;
    LAYER V1 ;
      RECT 8064 2712 8096 2744 ;
    LAYER V1 ;
      RECT 8064 2840 8096 2872 ;
    LAYER V1 ;
      RECT 8064 2968 8096 3000 ;
    LAYER V1 ;
      RECT 8064 3096 8096 3128 ;
    LAYER V1 ;
      RECT 8064 3224 8096 3256 ;
    LAYER V1 ;
      RECT 8064 3352 8096 3384 ;
    LAYER V1 ;
      RECT 8064 3480 8096 3512 ;
    LAYER V1 ;
      RECT 8064 3608 8096 3640 ;
    LAYER V1 ;
      RECT 8064 3736 8096 3768 ;
    LAYER V1 ;
      RECT 8064 3864 8096 3896 ;
    LAYER V1 ;
      RECT 8064 3992 8096 4024 ;
    LAYER V1 ;
      RECT 8064 4120 8096 4152 ;
    LAYER V1 ;
      RECT 8064 4248 8096 4280 ;
    LAYER V1 ;
      RECT 8064 4376 8096 4408 ;
    LAYER V1 ;
      RECT 8064 4504 8096 4536 ;
    LAYER V1 ;
      RECT 8064 4632 8096 4664 ;
    LAYER V1 ;
      RECT 8064 4760 8096 4792 ;
    LAYER V1 ;
      RECT 8064 4888 8096 4920 ;
    LAYER V1 ;
      RECT 8064 5016 8096 5048 ;
    LAYER V1 ;
      RECT 8064 5144 8096 5176 ;
    LAYER V1 ;
      RECT 8064 5272 8096 5304 ;
    LAYER V1 ;
      RECT 8064 5400 8096 5432 ;
    LAYER V1 ;
      RECT 8064 5528 8096 5560 ;
    LAYER V1 ;
      RECT 8064 5656 8096 5688 ;
    LAYER V1 ;
      RECT 8064 5784 8096 5816 ;
    LAYER V1 ;
      RECT 8064 5912 8096 5944 ;
    LAYER V1 ;
      RECT 8064 6040 8096 6072 ;
    LAYER V1 ;
      RECT 8064 6168 8096 6200 ;
    LAYER V1 ;
      RECT 8064 6296 8096 6328 ;
    LAYER V1 ;
      RECT 8064 6424 8096 6456 ;
    LAYER V1 ;
      RECT 8064 6552 8096 6584 ;
    LAYER V1 ;
      RECT 8064 6680 8096 6712 ;
    LAYER V1 ;
      RECT 8064 6808 8096 6840 ;
    LAYER V1 ;
      RECT 8064 6936 8096 6968 ;
    LAYER V1 ;
      RECT 8064 7064 8096 7096 ;
    LAYER V1 ;
      RECT 8064 7192 8096 7224 ;
    LAYER V1 ;
      RECT 8064 7320 8096 7352 ;
    LAYER V1 ;
      RECT 8064 7448 8096 7480 ;
    LAYER V1 ;
      RECT 8064 7576 8096 7608 ;
    LAYER V1 ;
      RECT 8064 7704 8096 7736 ;
    LAYER V1 ;
      RECT 8064 7832 8096 7864 ;
    LAYER M3 ;
      RECT 304 132 336 8016 ;
    LAYER M3 ;
      RECT 368 132 400 8016 ;
    LAYER M3 ;
      RECT 432 132 464 8016 ;
    LAYER M3 ;
      RECT 496 132 528 8016 ;
    LAYER M3 ;
      RECT 560 132 592 8016 ;
    LAYER M3 ;
      RECT 624 132 656 8016 ;
    LAYER M3 ;
      RECT 688 132 720 8016 ;
    LAYER M3 ;
      RECT 752 132 784 8016 ;
    LAYER M3 ;
      RECT 816 132 848 8016 ;
    LAYER M3 ;
      RECT 880 132 912 8016 ;
    LAYER M3 ;
      RECT 944 132 976 8016 ;
    LAYER M3 ;
      RECT 1008 132 1040 8016 ;
    LAYER M3 ;
      RECT 1072 132 1104 8016 ;
    LAYER M3 ;
      RECT 1136 132 1168 8016 ;
    LAYER M3 ;
      RECT 1200 132 1232 8016 ;
    LAYER M3 ;
      RECT 1264 132 1296 8016 ;
    LAYER M3 ;
      RECT 1328 132 1360 8016 ;
    LAYER M3 ;
      RECT 1392 132 1424 8016 ;
    LAYER M3 ;
      RECT 1456 132 1488 8016 ;
    LAYER M3 ;
      RECT 1520 132 1552 8016 ;
    LAYER M3 ;
      RECT 1584 132 1616 8016 ;
    LAYER M3 ;
      RECT 1648 132 1680 8016 ;
    LAYER M3 ;
      RECT 1712 132 1744 8016 ;
    LAYER M3 ;
      RECT 1776 132 1808 8016 ;
    LAYER M3 ;
      RECT 1840 132 1872 8016 ;
    LAYER M3 ;
      RECT 1904 132 1936 8016 ;
    LAYER M3 ;
      RECT 1968 132 2000 8016 ;
    LAYER M3 ;
      RECT 2032 132 2064 8016 ;
    LAYER M3 ;
      RECT 2096 132 2128 8016 ;
    LAYER M3 ;
      RECT 2160 132 2192 8016 ;
    LAYER M3 ;
      RECT 2224 132 2256 8016 ;
    LAYER M3 ;
      RECT 2288 132 2320 8016 ;
    LAYER M3 ;
      RECT 2352 132 2384 8016 ;
    LAYER M3 ;
      RECT 2416 132 2448 8016 ;
    LAYER M3 ;
      RECT 2480 132 2512 8016 ;
    LAYER M3 ;
      RECT 2544 132 2576 8016 ;
    LAYER M3 ;
      RECT 2608 132 2640 8016 ;
    LAYER M3 ;
      RECT 2672 132 2704 8016 ;
    LAYER M3 ;
      RECT 2736 132 2768 8016 ;
    LAYER M3 ;
      RECT 2800 132 2832 8016 ;
    LAYER M3 ;
      RECT 2864 132 2896 8016 ;
    LAYER M3 ;
      RECT 2928 132 2960 8016 ;
    LAYER M3 ;
      RECT 2992 132 3024 8016 ;
    LAYER M3 ;
      RECT 3056 132 3088 8016 ;
    LAYER M3 ;
      RECT 3120 132 3152 8016 ;
    LAYER M3 ;
      RECT 3184 132 3216 8016 ;
    LAYER M3 ;
      RECT 3248 132 3280 8016 ;
    LAYER M3 ;
      RECT 3312 132 3344 8016 ;
    LAYER M3 ;
      RECT 3376 132 3408 8016 ;
    LAYER M3 ;
      RECT 3440 132 3472 8016 ;
    LAYER M3 ;
      RECT 3504 132 3536 8016 ;
    LAYER M3 ;
      RECT 3568 132 3600 8016 ;
    LAYER M3 ;
      RECT 3632 132 3664 8016 ;
    LAYER M3 ;
      RECT 3696 132 3728 8016 ;
    LAYER M3 ;
      RECT 3760 132 3792 8016 ;
    LAYER M3 ;
      RECT 3824 132 3856 8016 ;
    LAYER M3 ;
      RECT 3888 132 3920 8016 ;
    LAYER M3 ;
      RECT 3952 132 3984 8016 ;
    LAYER M3 ;
      RECT 4016 132 4048 8016 ;
    LAYER M3 ;
      RECT 4080 132 4112 8016 ;
    LAYER M3 ;
      RECT 4144 132 4176 8016 ;
    LAYER M3 ;
      RECT 4208 132 4240 8016 ;
    LAYER M3 ;
      RECT 4272 132 4304 8016 ;
    LAYER M3 ;
      RECT 4336 132 4368 8016 ;
    LAYER M3 ;
      RECT 4400 132 4432 8016 ;
    LAYER M3 ;
      RECT 4464 132 4496 8016 ;
    LAYER M3 ;
      RECT 4528 132 4560 8016 ;
    LAYER M3 ;
      RECT 4592 132 4624 8016 ;
    LAYER M3 ;
      RECT 4656 132 4688 8016 ;
    LAYER M3 ;
      RECT 4720 132 4752 8016 ;
    LAYER M3 ;
      RECT 4784 132 4816 8016 ;
    LAYER M3 ;
      RECT 4848 132 4880 8016 ;
    LAYER M3 ;
      RECT 4912 132 4944 8016 ;
    LAYER M3 ;
      RECT 4976 132 5008 8016 ;
    LAYER M3 ;
      RECT 5040 132 5072 8016 ;
    LAYER M3 ;
      RECT 5104 132 5136 8016 ;
    LAYER M3 ;
      RECT 5168 132 5200 8016 ;
    LAYER M3 ;
      RECT 5232 132 5264 8016 ;
    LAYER M3 ;
      RECT 5296 132 5328 8016 ;
    LAYER M3 ;
      RECT 5360 132 5392 8016 ;
    LAYER M3 ;
      RECT 5424 132 5456 8016 ;
    LAYER M3 ;
      RECT 5488 132 5520 8016 ;
    LAYER M3 ;
      RECT 5552 132 5584 8016 ;
    LAYER M3 ;
      RECT 5616 132 5648 8016 ;
    LAYER M3 ;
      RECT 5680 132 5712 8016 ;
    LAYER M3 ;
      RECT 5744 132 5776 8016 ;
    LAYER M3 ;
      RECT 5808 132 5840 8016 ;
    LAYER M3 ;
      RECT 5872 132 5904 8016 ;
    LAYER M3 ;
      RECT 5936 132 5968 8016 ;
    LAYER M3 ;
      RECT 6000 132 6032 8016 ;
    LAYER M3 ;
      RECT 6064 132 6096 8016 ;
    LAYER M3 ;
      RECT 6128 132 6160 8016 ;
    LAYER M3 ;
      RECT 6192 132 6224 8016 ;
    LAYER M3 ;
      RECT 6256 132 6288 8016 ;
    LAYER M3 ;
      RECT 6320 132 6352 8016 ;
    LAYER M3 ;
      RECT 6384 132 6416 8016 ;
    LAYER M3 ;
      RECT 6448 132 6480 8016 ;
    LAYER M3 ;
      RECT 6512 132 6544 8016 ;
    LAYER M3 ;
      RECT 6576 132 6608 8016 ;
    LAYER M3 ;
      RECT 6640 132 6672 8016 ;
    LAYER M3 ;
      RECT 6704 132 6736 8016 ;
    LAYER M3 ;
      RECT 6768 132 6800 8016 ;
    LAYER M3 ;
      RECT 6832 132 6864 8016 ;
    LAYER M3 ;
      RECT 6896 132 6928 8016 ;
    LAYER M3 ;
      RECT 6960 132 6992 8016 ;
    LAYER M3 ;
      RECT 7024 132 7056 8016 ;
    LAYER M3 ;
      RECT 7088 132 7120 8016 ;
    LAYER M3 ;
      RECT 7152 132 7184 8016 ;
    LAYER M3 ;
      RECT 7216 132 7248 8016 ;
    LAYER M3 ;
      RECT 7280 132 7312 8016 ;
    LAYER M3 ;
      RECT 7344 132 7376 8016 ;
    LAYER M3 ;
      RECT 7408 132 7440 8016 ;
    LAYER M3 ;
      RECT 7472 132 7504 8016 ;
    LAYER M3 ;
      RECT 7536 132 7568 8016 ;
    LAYER M3 ;
      RECT 7600 132 7632 8016 ;
    LAYER M3 ;
      RECT 7664 132 7696 8016 ;
    LAYER M3 ;
      RECT 7728 132 7760 8016 ;
    LAYER M3 ;
      RECT 7792 132 7824 8016 ;
    LAYER M3 ;
      RECT 7856 132 7888 8016 ;
    LAYER M3 ;
      RECT 7920 132 7952 8016 ;
    LAYER M3 ;
      RECT 7984 132 8016 8016 ;
    LAYER M3 ;
      RECT 8060 132 8100 8016 ;
    LAYER V2 ;
      RECT 304 216 336 248 ;
    LAYER V2 ;
      RECT 304 344 336 376 ;
    LAYER V2 ;
      RECT 304 472 336 504 ;
    LAYER V2 ;
      RECT 304 600 336 632 ;
    LAYER V2 ;
      RECT 304 728 336 760 ;
    LAYER V2 ;
      RECT 304 856 336 888 ;
    LAYER V2 ;
      RECT 304 984 336 1016 ;
    LAYER V2 ;
      RECT 304 1112 336 1144 ;
    LAYER V2 ;
      RECT 304 1240 336 1272 ;
    LAYER V2 ;
      RECT 304 1368 336 1400 ;
    LAYER V2 ;
      RECT 304 1496 336 1528 ;
    LAYER V2 ;
      RECT 304 1624 336 1656 ;
    LAYER V2 ;
      RECT 304 1752 336 1784 ;
    LAYER V2 ;
      RECT 304 1880 336 1912 ;
    LAYER V2 ;
      RECT 304 2008 336 2040 ;
    LAYER V2 ;
      RECT 304 2136 336 2168 ;
    LAYER V2 ;
      RECT 304 2264 336 2296 ;
    LAYER V2 ;
      RECT 304 2392 336 2424 ;
    LAYER V2 ;
      RECT 304 2520 336 2552 ;
    LAYER V2 ;
      RECT 304 2648 336 2680 ;
    LAYER V2 ;
      RECT 304 2776 336 2808 ;
    LAYER V2 ;
      RECT 304 2904 336 2936 ;
    LAYER V2 ;
      RECT 304 3032 336 3064 ;
    LAYER V2 ;
      RECT 304 3160 336 3192 ;
    LAYER V2 ;
      RECT 304 3288 336 3320 ;
    LAYER V2 ;
      RECT 304 3416 336 3448 ;
    LAYER V2 ;
      RECT 304 3544 336 3576 ;
    LAYER V2 ;
      RECT 304 3672 336 3704 ;
    LAYER V2 ;
      RECT 304 3800 336 3832 ;
    LAYER V2 ;
      RECT 304 3928 336 3960 ;
    LAYER V2 ;
      RECT 304 4056 336 4088 ;
    LAYER V2 ;
      RECT 304 4184 336 4216 ;
    LAYER V2 ;
      RECT 304 4312 336 4344 ;
    LAYER V2 ;
      RECT 304 4440 336 4472 ;
    LAYER V2 ;
      RECT 304 4568 336 4600 ;
    LAYER V2 ;
      RECT 304 4696 336 4728 ;
    LAYER V2 ;
      RECT 304 4824 336 4856 ;
    LAYER V2 ;
      RECT 304 4952 336 4984 ;
    LAYER V2 ;
      RECT 304 5080 336 5112 ;
    LAYER V2 ;
      RECT 304 5208 336 5240 ;
    LAYER V2 ;
      RECT 304 5336 336 5368 ;
    LAYER V2 ;
      RECT 304 5464 336 5496 ;
    LAYER V2 ;
      RECT 304 5592 336 5624 ;
    LAYER V2 ;
      RECT 304 5720 336 5752 ;
    LAYER V2 ;
      RECT 304 5848 336 5880 ;
    LAYER V2 ;
      RECT 304 5976 336 6008 ;
    LAYER V2 ;
      RECT 304 6104 336 6136 ;
    LAYER V2 ;
      RECT 304 6232 336 6264 ;
    LAYER V2 ;
      RECT 304 6360 336 6392 ;
    LAYER V2 ;
      RECT 304 6488 336 6520 ;
    LAYER V2 ;
      RECT 304 6616 336 6648 ;
    LAYER V2 ;
      RECT 304 6744 336 6776 ;
    LAYER V2 ;
      RECT 304 6872 336 6904 ;
    LAYER V2 ;
      RECT 304 7000 336 7032 ;
    LAYER V2 ;
      RECT 304 7128 336 7160 ;
    LAYER V2 ;
      RECT 304 7256 336 7288 ;
    LAYER V2 ;
      RECT 304 7384 336 7416 ;
    LAYER V2 ;
      RECT 304 7512 336 7544 ;
    LAYER V2 ;
      RECT 304 7640 336 7672 ;
    LAYER V2 ;
      RECT 304 7768 336 7800 ;
    LAYER V2 ;
      RECT 304 7964 336 7996 ;
    LAYER V2 ;
      RECT 368 152 400 184 ;
    LAYER V2 ;
      RECT 432 7964 464 7996 ;
    LAYER V2 ;
      RECT 496 152 528 184 ;
    LAYER V2 ;
      RECT 560 7964 592 7996 ;
    LAYER V2 ;
      RECT 624 152 656 184 ;
    LAYER V2 ;
      RECT 688 7964 720 7996 ;
    LAYER V2 ;
      RECT 752 152 784 184 ;
    LAYER V2 ;
      RECT 816 7964 848 7996 ;
    LAYER V2 ;
      RECT 880 152 912 184 ;
    LAYER V2 ;
      RECT 944 7964 976 7996 ;
    LAYER V2 ;
      RECT 1008 152 1040 184 ;
    LAYER V2 ;
      RECT 1072 7964 1104 7996 ;
    LAYER V2 ;
      RECT 1136 152 1168 184 ;
    LAYER V2 ;
      RECT 1200 7964 1232 7996 ;
    LAYER V2 ;
      RECT 1264 152 1296 184 ;
    LAYER V2 ;
      RECT 1328 7964 1360 7996 ;
    LAYER V2 ;
      RECT 1392 152 1424 184 ;
    LAYER V2 ;
      RECT 1456 7964 1488 7996 ;
    LAYER V2 ;
      RECT 1520 152 1552 184 ;
    LAYER V2 ;
      RECT 1584 7964 1616 7996 ;
    LAYER V2 ;
      RECT 1648 152 1680 184 ;
    LAYER V2 ;
      RECT 1712 7964 1744 7996 ;
    LAYER V2 ;
      RECT 1776 152 1808 184 ;
    LAYER V2 ;
      RECT 1840 7964 1872 7996 ;
    LAYER V2 ;
      RECT 1904 152 1936 184 ;
    LAYER V2 ;
      RECT 1968 7964 2000 7996 ;
    LAYER V2 ;
      RECT 2032 152 2064 184 ;
    LAYER V2 ;
      RECT 2096 7964 2128 7996 ;
    LAYER V2 ;
      RECT 2160 152 2192 184 ;
    LAYER V2 ;
      RECT 2224 7964 2256 7996 ;
    LAYER V2 ;
      RECT 2288 152 2320 184 ;
    LAYER V2 ;
      RECT 2352 7964 2384 7996 ;
    LAYER V2 ;
      RECT 2416 152 2448 184 ;
    LAYER V2 ;
      RECT 2480 7964 2512 7996 ;
    LAYER V2 ;
      RECT 2544 152 2576 184 ;
    LAYER V2 ;
      RECT 2608 7964 2640 7996 ;
    LAYER V2 ;
      RECT 2672 152 2704 184 ;
    LAYER V2 ;
      RECT 2736 7964 2768 7996 ;
    LAYER V2 ;
      RECT 2800 152 2832 184 ;
    LAYER V2 ;
      RECT 2864 7964 2896 7996 ;
    LAYER V2 ;
      RECT 2928 152 2960 184 ;
    LAYER V2 ;
      RECT 2992 7964 3024 7996 ;
    LAYER V2 ;
      RECT 3056 152 3088 184 ;
    LAYER V2 ;
      RECT 3120 7964 3152 7996 ;
    LAYER V2 ;
      RECT 3184 152 3216 184 ;
    LAYER V2 ;
      RECT 3248 7964 3280 7996 ;
    LAYER V2 ;
      RECT 3312 152 3344 184 ;
    LAYER V2 ;
      RECT 3376 7964 3408 7996 ;
    LAYER V2 ;
      RECT 3440 152 3472 184 ;
    LAYER V2 ;
      RECT 3504 7964 3536 7996 ;
    LAYER V2 ;
      RECT 3568 152 3600 184 ;
    LAYER V2 ;
      RECT 3632 7964 3664 7996 ;
    LAYER V2 ;
      RECT 3696 152 3728 184 ;
    LAYER V2 ;
      RECT 3760 7964 3792 7996 ;
    LAYER V2 ;
      RECT 3824 152 3856 184 ;
    LAYER V2 ;
      RECT 3888 7964 3920 7996 ;
    LAYER V2 ;
      RECT 3952 152 3984 184 ;
    LAYER V2 ;
      RECT 4016 7964 4048 7996 ;
    LAYER V2 ;
      RECT 4080 152 4112 184 ;
    LAYER V2 ;
      RECT 4144 7964 4176 7996 ;
    LAYER V2 ;
      RECT 4208 152 4240 184 ;
    LAYER V2 ;
      RECT 4272 7964 4304 7996 ;
    LAYER V2 ;
      RECT 4336 152 4368 184 ;
    LAYER V2 ;
      RECT 4400 7964 4432 7996 ;
    LAYER V2 ;
      RECT 4464 152 4496 184 ;
    LAYER V2 ;
      RECT 4528 7964 4560 7996 ;
    LAYER V2 ;
      RECT 4592 152 4624 184 ;
    LAYER V2 ;
      RECT 4656 7964 4688 7996 ;
    LAYER V2 ;
      RECT 4720 152 4752 184 ;
    LAYER V2 ;
      RECT 4784 7964 4816 7996 ;
    LAYER V2 ;
      RECT 4848 152 4880 184 ;
    LAYER V2 ;
      RECT 4912 7964 4944 7996 ;
    LAYER V2 ;
      RECT 4976 152 5008 184 ;
    LAYER V2 ;
      RECT 5040 7964 5072 7996 ;
    LAYER V2 ;
      RECT 5104 152 5136 184 ;
    LAYER V2 ;
      RECT 5168 7964 5200 7996 ;
    LAYER V2 ;
      RECT 5232 152 5264 184 ;
    LAYER V2 ;
      RECT 5296 7964 5328 7996 ;
    LAYER V2 ;
      RECT 5360 152 5392 184 ;
    LAYER V2 ;
      RECT 5424 7964 5456 7996 ;
    LAYER V2 ;
      RECT 5488 152 5520 184 ;
    LAYER V2 ;
      RECT 5552 7964 5584 7996 ;
    LAYER V2 ;
      RECT 5616 152 5648 184 ;
    LAYER V2 ;
      RECT 5680 7964 5712 7996 ;
    LAYER V2 ;
      RECT 5744 152 5776 184 ;
    LAYER V2 ;
      RECT 5808 7964 5840 7996 ;
    LAYER V2 ;
      RECT 5872 152 5904 184 ;
    LAYER V2 ;
      RECT 5936 7964 5968 7996 ;
    LAYER V2 ;
      RECT 6000 152 6032 184 ;
    LAYER V2 ;
      RECT 6064 7964 6096 7996 ;
    LAYER V2 ;
      RECT 6128 152 6160 184 ;
    LAYER V2 ;
      RECT 6192 7964 6224 7996 ;
    LAYER V2 ;
      RECT 6256 152 6288 184 ;
    LAYER V2 ;
      RECT 6320 7964 6352 7996 ;
    LAYER V2 ;
      RECT 6384 152 6416 184 ;
    LAYER V2 ;
      RECT 6448 7964 6480 7996 ;
    LAYER V2 ;
      RECT 6512 152 6544 184 ;
    LAYER V2 ;
      RECT 6576 7964 6608 7996 ;
    LAYER V2 ;
      RECT 6640 152 6672 184 ;
    LAYER V2 ;
      RECT 6704 7964 6736 7996 ;
    LAYER V2 ;
      RECT 6768 152 6800 184 ;
    LAYER V2 ;
      RECT 6832 7964 6864 7996 ;
    LAYER V2 ;
      RECT 6896 152 6928 184 ;
    LAYER V2 ;
      RECT 6960 7964 6992 7996 ;
    LAYER V2 ;
      RECT 7024 152 7056 184 ;
    LAYER V2 ;
      RECT 7088 7964 7120 7996 ;
    LAYER V2 ;
      RECT 7152 152 7184 184 ;
    LAYER V2 ;
      RECT 7216 7964 7248 7996 ;
    LAYER V2 ;
      RECT 7280 152 7312 184 ;
    LAYER V2 ;
      RECT 7344 7964 7376 7996 ;
    LAYER V2 ;
      RECT 7408 152 7440 184 ;
    LAYER V2 ;
      RECT 7472 7964 7504 7996 ;
    LAYER V2 ;
      RECT 7536 152 7568 184 ;
    LAYER V2 ;
      RECT 7600 7964 7632 7996 ;
    LAYER V2 ;
      RECT 7664 152 7696 184 ;
    LAYER V2 ;
      RECT 7728 7964 7760 7996 ;
    LAYER V2 ;
      RECT 7792 152 7824 184 ;
    LAYER V2 ;
      RECT 7856 7964 7888 7996 ;
    LAYER V2 ;
      RECT 7920 152 7952 184 ;
    LAYER V2 ;
      RECT 7984 7964 8016 7996 ;
    LAYER V2 ;
      RECT 8064 152 8096 184 ;
    LAYER V2 ;
      RECT 8064 280 8096 312 ;
    LAYER V2 ;
      RECT 8064 408 8096 440 ;
    LAYER V2 ;
      RECT 8064 536 8096 568 ;
    LAYER V2 ;
      RECT 8064 664 8096 696 ;
    LAYER V2 ;
      RECT 8064 792 8096 824 ;
    LAYER V2 ;
      RECT 8064 920 8096 952 ;
    LAYER V2 ;
      RECT 8064 1048 8096 1080 ;
    LAYER V2 ;
      RECT 8064 1176 8096 1208 ;
    LAYER V2 ;
      RECT 8064 1304 8096 1336 ;
    LAYER V2 ;
      RECT 8064 1432 8096 1464 ;
    LAYER V2 ;
      RECT 8064 1560 8096 1592 ;
    LAYER V2 ;
      RECT 8064 1688 8096 1720 ;
    LAYER V2 ;
      RECT 8064 1816 8096 1848 ;
    LAYER V2 ;
      RECT 8064 1944 8096 1976 ;
    LAYER V2 ;
      RECT 8064 2072 8096 2104 ;
    LAYER V2 ;
      RECT 8064 2200 8096 2232 ;
    LAYER V2 ;
      RECT 8064 2328 8096 2360 ;
    LAYER V2 ;
      RECT 8064 2456 8096 2488 ;
    LAYER V2 ;
      RECT 8064 2584 8096 2616 ;
    LAYER V2 ;
      RECT 8064 2712 8096 2744 ;
    LAYER V2 ;
      RECT 8064 2840 8096 2872 ;
    LAYER V2 ;
      RECT 8064 2968 8096 3000 ;
    LAYER V2 ;
      RECT 8064 3096 8096 3128 ;
    LAYER V2 ;
      RECT 8064 3224 8096 3256 ;
    LAYER V2 ;
      RECT 8064 3352 8096 3384 ;
    LAYER V2 ;
      RECT 8064 3480 8096 3512 ;
    LAYER V2 ;
      RECT 8064 3608 8096 3640 ;
    LAYER V2 ;
      RECT 8064 3736 8096 3768 ;
    LAYER V2 ;
      RECT 8064 3864 8096 3896 ;
    LAYER V2 ;
      RECT 8064 3992 8096 4024 ;
    LAYER V2 ;
      RECT 8064 4120 8096 4152 ;
    LAYER V2 ;
      RECT 8064 4248 8096 4280 ;
    LAYER V2 ;
      RECT 8064 4376 8096 4408 ;
    LAYER V2 ;
      RECT 8064 4504 8096 4536 ;
    LAYER V2 ;
      RECT 8064 4632 8096 4664 ;
    LAYER V2 ;
      RECT 8064 4760 8096 4792 ;
    LAYER V2 ;
      RECT 8064 4888 8096 4920 ;
    LAYER V2 ;
      RECT 8064 5016 8096 5048 ;
    LAYER V2 ;
      RECT 8064 5144 8096 5176 ;
    LAYER V2 ;
      RECT 8064 5272 8096 5304 ;
    LAYER V2 ;
      RECT 8064 5400 8096 5432 ;
    LAYER V2 ;
      RECT 8064 5528 8096 5560 ;
    LAYER V2 ;
      RECT 8064 5656 8096 5688 ;
    LAYER V2 ;
      RECT 8064 5784 8096 5816 ;
    LAYER V2 ;
      RECT 8064 5912 8096 5944 ;
    LAYER V2 ;
      RECT 8064 6040 8096 6072 ;
    LAYER V2 ;
      RECT 8064 6168 8096 6200 ;
    LAYER V2 ;
      RECT 8064 6296 8096 6328 ;
    LAYER V2 ;
      RECT 8064 6424 8096 6456 ;
    LAYER V2 ;
      RECT 8064 6552 8096 6584 ;
    LAYER V2 ;
      RECT 8064 6680 8096 6712 ;
    LAYER V2 ;
      RECT 8064 6808 8096 6840 ;
    LAYER V2 ;
      RECT 8064 6936 8096 6968 ;
    LAYER V2 ;
      RECT 8064 7064 8096 7096 ;
    LAYER V2 ;
      RECT 8064 7192 8096 7224 ;
    LAYER V2 ;
      RECT 8064 7320 8096 7352 ;
    LAYER V2 ;
      RECT 8064 7448 8096 7480 ;
    LAYER V2 ;
      RECT 8064 7576 8096 7608 ;
    LAYER V2 ;
      RECT 8064 7704 8096 7736 ;
    LAYER V2 ;
      RECT 8064 7832 8096 7864 ;
  END
END CAP_12F
MACRO CMC_NMOS_B_97926084_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CMC_NMOS_B_97926084_X1_Y1 0 0 ;
  SIZE 800 BY 2352 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 1748 516 1780 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124 68 356 100 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 152 516 184 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 908 516 940 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204 236 596 268 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1644 336 1884 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 464 48 496 792 ;
    LAYER M1 ;
      RECT 464 888 496 1128 ;
    LAYER M1 ;
      RECT 464 1644 496 1884 ;
    LAYER M1 ;
      RECT 544 48 576 792 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1748 336 1780 ;
    LAYER V1 ;
      RECT 464 152 496 184 ;
    LAYER V1 ;
      RECT 464 908 496 940 ;
    LAYER V1 ;
      RECT 464 1748 496 1780 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 544 236 576 268 ;
    LAYER V0 ;
      RECT 304 461 336 493 ;
    LAYER V0 ;
      RECT 304 545 336 577 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1748 336 1780 ;
    LAYER V0 ;
      RECT 224 461 256 493 ;
    LAYER V0 ;
      RECT 224 545 256 577 ;
    LAYER V0 ;
      RECT 384 461 416 493 ;
    LAYER V0 ;
      RECT 384 461 416 493 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 464 461 496 493 ;
    LAYER V0 ;
      RECT 464 545 496 577 ;
    LAYER V0 ;
      RECT 464 908 496 940 ;
    LAYER V0 ;
      RECT 464 1748 496 1780 ;
    LAYER V0 ;
      RECT 544 461 576 493 ;
    LAYER V0 ;
      RECT 544 545 576 577 ;
  END
END CMC_NMOS_B_97926084_X1_Y1
MACRO CMC_S_NMOS_B_94218540_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CMC_S_NMOS_B_94218540_X1_Y1 0 0 ;
  SIZE 1280 BY 2352 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 1748 996 1780 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 68 516 100 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 764 152 996 184 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 908 996 940 ;
    END
  END G
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204 236 436 268 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 844 320 1076 352 ;
    END
  END SB
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1644 336 1884 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 944 48 976 792 ;
    LAYER M1 ;
      RECT 944 888 976 1128 ;
    LAYER M1 ;
      RECT 944 1644 976 1884 ;
    LAYER M1 ;
      RECT 864 48 896 792 ;
    LAYER M1 ;
      RECT 1024 48 1056 792 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1748 336 1780 ;
    LAYER V1 ;
      RECT 944 152 976 184 ;
    LAYER V1 ;
      RECT 944 908 976 940 ;
    LAYER V1 ;
      RECT 944 1748 976 1780 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 864 320 896 352 ;
    LAYER V1 ;
      RECT 1024 320 1056 352 ;
    LAYER V0 ;
      RECT 304 461 336 493 ;
    LAYER V0 ;
      RECT 304 545 336 577 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1748 336 1780 ;
    LAYER V0 ;
      RECT 224 461 256 493 ;
    LAYER V0 ;
      RECT 224 545 256 577 ;
    LAYER V0 ;
      RECT 384 461 416 493 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 944 461 976 493 ;
    LAYER V0 ;
      RECT 944 545 976 577 ;
    LAYER V0 ;
      RECT 944 908 976 940 ;
    LAYER V0 ;
      RECT 944 1748 976 1780 ;
    LAYER V0 ;
      RECT 864 461 896 493 ;
    LAYER V0 ;
      RECT 864 545 896 577 ;
    LAYER V0 ;
      RECT 1024 461 1056 493 ;
    LAYER V0 ;
      RECT 1024 545 1056 577 ;
  END
END CMC_S_NMOS_B_94218540_X1_Y1
MACRO CAP_2T_57809468
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CAP_2T_57809468 0 0 ;
  SIZE 6080 BY 5796 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44 5612 6036 5644 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44 152 6036 184 ;
    END
  END PLUS
  OBS
    LAYER M1 ;
      RECT 304 132 336 5664 ;
    LAYER M1 ;
      RECT 368 132 400 5664 ;
    LAYER M1 ;
      RECT 432 132 464 5664 ;
    LAYER M1 ;
      RECT 496 132 528 5664 ;
    LAYER M1 ;
      RECT 560 132 592 5664 ;
    LAYER M1 ;
      RECT 624 132 656 5664 ;
    LAYER M1 ;
      RECT 688 132 720 5664 ;
    LAYER M1 ;
      RECT 752 132 784 5664 ;
    LAYER M1 ;
      RECT 816 132 848 5664 ;
    LAYER M1 ;
      RECT 880 132 912 5664 ;
    LAYER M1 ;
      RECT 944 132 976 5664 ;
    LAYER M1 ;
      RECT 1008 132 1040 5664 ;
    LAYER M1 ;
      RECT 1072 132 1104 5664 ;
    LAYER M1 ;
      RECT 1136 132 1168 5664 ;
    LAYER M1 ;
      RECT 1200 132 1232 5664 ;
    LAYER M1 ;
      RECT 1264 132 1296 5664 ;
    LAYER M1 ;
      RECT 1328 132 1360 5664 ;
    LAYER M1 ;
      RECT 1392 132 1424 5664 ;
    LAYER M1 ;
      RECT 1456 132 1488 5664 ;
    LAYER M1 ;
      RECT 1520 132 1552 5664 ;
    LAYER M1 ;
      RECT 1584 132 1616 5664 ;
    LAYER M1 ;
      RECT 1648 132 1680 5664 ;
    LAYER M1 ;
      RECT 1712 132 1744 5664 ;
    LAYER M1 ;
      RECT 1776 132 1808 5664 ;
    LAYER M1 ;
      RECT 1840 132 1872 5664 ;
    LAYER M1 ;
      RECT 1904 132 1936 5664 ;
    LAYER M1 ;
      RECT 1968 132 2000 5664 ;
    LAYER M1 ;
      RECT 2032 132 2064 5664 ;
    LAYER M1 ;
      RECT 2096 132 2128 5664 ;
    LAYER M1 ;
      RECT 2160 132 2192 5664 ;
    LAYER M1 ;
      RECT 2224 132 2256 5664 ;
    LAYER M1 ;
      RECT 2288 132 2320 5664 ;
    LAYER M1 ;
      RECT 2352 132 2384 5664 ;
    LAYER M1 ;
      RECT 2416 132 2448 5664 ;
    LAYER M1 ;
      RECT 2480 132 2512 5664 ;
    LAYER M1 ;
      RECT 2544 132 2576 5664 ;
    LAYER M1 ;
      RECT 2608 132 2640 5664 ;
    LAYER M1 ;
      RECT 2672 132 2704 5664 ;
    LAYER M1 ;
      RECT 2736 132 2768 5664 ;
    LAYER M1 ;
      RECT 2800 132 2832 5664 ;
    LAYER M1 ;
      RECT 2864 132 2896 5664 ;
    LAYER M1 ;
      RECT 2928 132 2960 5664 ;
    LAYER M1 ;
      RECT 2992 132 3024 5664 ;
    LAYER M1 ;
      RECT 3056 132 3088 5664 ;
    LAYER M1 ;
      RECT 3120 132 3152 5664 ;
    LAYER M1 ;
      RECT 3184 132 3216 5664 ;
    LAYER M1 ;
      RECT 3248 132 3280 5664 ;
    LAYER M1 ;
      RECT 3312 132 3344 5664 ;
    LAYER M1 ;
      RECT 3376 132 3408 5664 ;
    LAYER M1 ;
      RECT 3440 132 3472 5664 ;
    LAYER M1 ;
      RECT 3504 132 3536 5664 ;
    LAYER M1 ;
      RECT 3568 132 3600 5664 ;
    LAYER M1 ;
      RECT 3632 132 3664 5664 ;
    LAYER M1 ;
      RECT 3696 132 3728 5664 ;
    LAYER M1 ;
      RECT 3760 132 3792 5664 ;
    LAYER M1 ;
      RECT 3824 132 3856 5664 ;
    LAYER M1 ;
      RECT 3888 132 3920 5664 ;
    LAYER M1 ;
      RECT 3952 132 3984 5664 ;
    LAYER M1 ;
      RECT 4016 132 4048 5664 ;
    LAYER M1 ;
      RECT 4080 132 4112 5664 ;
    LAYER M1 ;
      RECT 4144 132 4176 5664 ;
    LAYER M1 ;
      RECT 4208 132 4240 5664 ;
    LAYER M1 ;
      RECT 4272 132 4304 5664 ;
    LAYER M1 ;
      RECT 4336 132 4368 5664 ;
    LAYER M1 ;
      RECT 4400 132 4432 5664 ;
    LAYER M1 ;
      RECT 4464 132 4496 5664 ;
    LAYER M1 ;
      RECT 4528 132 4560 5664 ;
    LAYER M1 ;
      RECT 4592 132 4624 5664 ;
    LAYER M1 ;
      RECT 4656 132 4688 5664 ;
    LAYER M1 ;
      RECT 4720 132 4752 5664 ;
    LAYER M1 ;
      RECT 4784 132 4816 5664 ;
    LAYER M1 ;
      RECT 4848 132 4880 5664 ;
    LAYER M1 ;
      RECT 4912 132 4944 5664 ;
    LAYER M1 ;
      RECT 4976 132 5008 5664 ;
    LAYER M1 ;
      RECT 5040 132 5072 5664 ;
    LAYER M1 ;
      RECT 5104 132 5136 5664 ;
    LAYER M1 ;
      RECT 5168 132 5200 5664 ;
    LAYER M1 ;
      RECT 5232 132 5264 5664 ;
    LAYER M1 ;
      RECT 5296 132 5328 5664 ;
    LAYER M1 ;
      RECT 5360 132 5392 5664 ;
    LAYER M1 ;
      RECT 5424 132 5456 5664 ;
    LAYER M1 ;
      RECT 5488 132 5520 5664 ;
    LAYER M1 ;
      RECT 5552 132 5584 5664 ;
    LAYER M1 ;
      RECT 5616 132 5648 5664 ;
    LAYER M1 ;
      RECT 5680 132 5712 5664 ;
    LAYER M1 ;
      RECT 5744 132 5776 5664 ;
    LAYER M2 ;
      RECT 284 216 5796 248 ;
    LAYER M2 ;
      RECT 284 280 5796 312 ;
    LAYER M2 ;
      RECT 284 344 5796 376 ;
    LAYER M2 ;
      RECT 284 408 5796 440 ;
    LAYER M2 ;
      RECT 284 472 5796 504 ;
    LAYER M2 ;
      RECT 284 536 5796 568 ;
    LAYER M2 ;
      RECT 284 600 5796 632 ;
    LAYER M2 ;
      RECT 284 664 5796 696 ;
    LAYER M2 ;
      RECT 284 728 5796 760 ;
    LAYER M2 ;
      RECT 284 792 5796 824 ;
    LAYER M2 ;
      RECT 284 856 5796 888 ;
    LAYER M2 ;
      RECT 284 920 5796 952 ;
    LAYER M2 ;
      RECT 284 984 5796 1016 ;
    LAYER M2 ;
      RECT 284 1048 5796 1080 ;
    LAYER M2 ;
      RECT 284 1112 5796 1144 ;
    LAYER M2 ;
      RECT 284 1176 5796 1208 ;
    LAYER M2 ;
      RECT 284 1240 5796 1272 ;
    LAYER M2 ;
      RECT 284 1304 5796 1336 ;
    LAYER M2 ;
      RECT 284 1368 5796 1400 ;
    LAYER M2 ;
      RECT 284 1432 5796 1464 ;
    LAYER M2 ;
      RECT 284 1496 5796 1528 ;
    LAYER M2 ;
      RECT 284 1560 5796 1592 ;
    LAYER M2 ;
      RECT 284 1624 5796 1656 ;
    LAYER M2 ;
      RECT 284 1688 5796 1720 ;
    LAYER M2 ;
      RECT 284 1752 5796 1784 ;
    LAYER M2 ;
      RECT 284 1816 5796 1848 ;
    LAYER M2 ;
      RECT 284 1880 5796 1912 ;
    LAYER M2 ;
      RECT 284 1944 5796 1976 ;
    LAYER M2 ;
      RECT 284 2008 5796 2040 ;
    LAYER M2 ;
      RECT 284 2072 5796 2104 ;
    LAYER M2 ;
      RECT 284 2136 5796 2168 ;
    LAYER M2 ;
      RECT 284 2200 5796 2232 ;
    LAYER M2 ;
      RECT 284 2264 5796 2296 ;
    LAYER M2 ;
      RECT 284 2328 5796 2360 ;
    LAYER M2 ;
      RECT 284 2392 5796 2424 ;
    LAYER M2 ;
      RECT 284 2456 5796 2488 ;
    LAYER M2 ;
      RECT 284 2520 5796 2552 ;
    LAYER M2 ;
      RECT 284 2584 5796 2616 ;
    LAYER M2 ;
      RECT 284 2648 5796 2680 ;
    LAYER M2 ;
      RECT 284 2712 5796 2744 ;
    LAYER M2 ;
      RECT 284 2776 5796 2808 ;
    LAYER M2 ;
      RECT 284 2840 5796 2872 ;
    LAYER M2 ;
      RECT 284 2904 5796 2936 ;
    LAYER M2 ;
      RECT 284 2968 5796 3000 ;
    LAYER M2 ;
      RECT 284 3032 5796 3064 ;
    LAYER M2 ;
      RECT 284 3096 5796 3128 ;
    LAYER M2 ;
      RECT 284 3160 5796 3192 ;
    LAYER M2 ;
      RECT 284 3224 5796 3256 ;
    LAYER M2 ;
      RECT 284 3288 5796 3320 ;
    LAYER M2 ;
      RECT 284 3352 5796 3384 ;
    LAYER M2 ;
      RECT 284 3416 5796 3448 ;
    LAYER M2 ;
      RECT 284 3480 5796 3512 ;
    LAYER M2 ;
      RECT 284 3544 5796 3576 ;
    LAYER M2 ;
      RECT 284 3608 5796 3640 ;
    LAYER M2 ;
      RECT 284 3672 5796 3704 ;
    LAYER M2 ;
      RECT 284 3736 5796 3768 ;
    LAYER M2 ;
      RECT 284 3800 5796 3832 ;
    LAYER M2 ;
      RECT 284 3864 5796 3896 ;
    LAYER M2 ;
      RECT 284 3928 5796 3960 ;
    LAYER M2 ;
      RECT 284 3992 5796 4024 ;
    LAYER M2 ;
      RECT 284 4056 5796 4088 ;
    LAYER M2 ;
      RECT 284 4120 5796 4152 ;
    LAYER M2 ;
      RECT 284 4184 5796 4216 ;
    LAYER M2 ;
      RECT 284 4248 5796 4280 ;
    LAYER M2 ;
      RECT 284 4312 5796 4344 ;
    LAYER M2 ;
      RECT 284 4376 5796 4408 ;
    LAYER M2 ;
      RECT 284 4440 5796 4472 ;
    LAYER M2 ;
      RECT 284 4504 5796 4536 ;
    LAYER M2 ;
      RECT 284 4568 5796 4600 ;
    LAYER M2 ;
      RECT 284 4632 5796 4664 ;
    LAYER M2 ;
      RECT 284 4696 5796 4728 ;
    LAYER M2 ;
      RECT 284 4760 5796 4792 ;
    LAYER M2 ;
      RECT 284 4824 5796 4856 ;
    LAYER M2 ;
      RECT 284 4888 5796 4920 ;
    LAYER M2 ;
      RECT 284 4952 5796 4984 ;
    LAYER M2 ;
      RECT 284 5016 5796 5048 ;
    LAYER M2 ;
      RECT 284 5080 5796 5112 ;
    LAYER M2 ;
      RECT 284 5144 5796 5176 ;
    LAYER M2 ;
      RECT 284 5208 5796 5240 ;
    LAYER M2 ;
      RECT 284 5272 5796 5304 ;
    LAYER M2 ;
      RECT 284 5336 5796 5368 ;
    LAYER M2 ;
      RECT 284 5400 5796 5432 ;
    LAYER M2 ;
      RECT 284 5464 5796 5496 ;
    LAYER M2 ;
      RECT 284 5528 5796 5560 ;
    LAYER V1 ;
      RECT 304 216 336 248 ;
    LAYER V1 ;
      RECT 304 344 336 376 ;
    LAYER V1 ;
      RECT 304 472 336 504 ;
    LAYER V1 ;
      RECT 304 600 336 632 ;
    LAYER V1 ;
      RECT 304 728 336 760 ;
    LAYER V1 ;
      RECT 304 856 336 888 ;
    LAYER V1 ;
      RECT 304 984 336 1016 ;
    LAYER V1 ;
      RECT 304 1112 336 1144 ;
    LAYER V1 ;
      RECT 304 1240 336 1272 ;
    LAYER V1 ;
      RECT 304 1368 336 1400 ;
    LAYER V1 ;
      RECT 304 1496 336 1528 ;
    LAYER V1 ;
      RECT 304 1624 336 1656 ;
    LAYER V1 ;
      RECT 304 1752 336 1784 ;
    LAYER V1 ;
      RECT 304 1880 336 1912 ;
    LAYER V1 ;
      RECT 304 2008 336 2040 ;
    LAYER V1 ;
      RECT 304 2136 336 2168 ;
    LAYER V1 ;
      RECT 304 2264 336 2296 ;
    LAYER V1 ;
      RECT 304 2392 336 2424 ;
    LAYER V1 ;
      RECT 304 2520 336 2552 ;
    LAYER V1 ;
      RECT 304 2648 336 2680 ;
    LAYER V1 ;
      RECT 304 2776 336 2808 ;
    LAYER V1 ;
      RECT 304 2904 336 2936 ;
    LAYER V1 ;
      RECT 304 3032 336 3064 ;
    LAYER V1 ;
      RECT 304 3160 336 3192 ;
    LAYER V1 ;
      RECT 304 3288 336 3320 ;
    LAYER V1 ;
      RECT 304 3416 336 3448 ;
    LAYER V1 ;
      RECT 304 3544 336 3576 ;
    LAYER V1 ;
      RECT 304 3672 336 3704 ;
    LAYER V1 ;
      RECT 304 3800 336 3832 ;
    LAYER V1 ;
      RECT 304 3928 336 3960 ;
    LAYER V1 ;
      RECT 304 4056 336 4088 ;
    LAYER V1 ;
      RECT 304 4184 336 4216 ;
    LAYER V1 ;
      RECT 304 4312 336 4344 ;
    LAYER V1 ;
      RECT 304 4440 336 4472 ;
    LAYER V1 ;
      RECT 304 4568 336 4600 ;
    LAYER V1 ;
      RECT 304 4696 336 4728 ;
    LAYER V1 ;
      RECT 304 4824 336 4856 ;
    LAYER V1 ;
      RECT 304 4952 336 4984 ;
    LAYER V1 ;
      RECT 304 5080 336 5112 ;
    LAYER V1 ;
      RECT 304 5208 336 5240 ;
    LAYER V1 ;
      RECT 304 5336 336 5368 ;
    LAYER V1 ;
      RECT 304 5464 336 5496 ;
    LAYER V1 ;
      RECT 304 5612 336 5644 ;
    LAYER V1 ;
      RECT 368 152 400 184 ;
    LAYER V1 ;
      RECT 432 5612 464 5644 ;
    LAYER V1 ;
      RECT 496 152 528 184 ;
    LAYER V1 ;
      RECT 560 5612 592 5644 ;
    LAYER V1 ;
      RECT 624 152 656 184 ;
    LAYER V1 ;
      RECT 688 5612 720 5644 ;
    LAYER V1 ;
      RECT 752 152 784 184 ;
    LAYER V1 ;
      RECT 816 5612 848 5644 ;
    LAYER V1 ;
      RECT 880 152 912 184 ;
    LAYER V1 ;
      RECT 944 5612 976 5644 ;
    LAYER V1 ;
      RECT 1008 152 1040 184 ;
    LAYER V1 ;
      RECT 1072 5612 1104 5644 ;
    LAYER V1 ;
      RECT 1136 152 1168 184 ;
    LAYER V1 ;
      RECT 1200 5612 1232 5644 ;
    LAYER V1 ;
      RECT 1264 152 1296 184 ;
    LAYER V1 ;
      RECT 1328 5612 1360 5644 ;
    LAYER V1 ;
      RECT 1392 152 1424 184 ;
    LAYER V1 ;
      RECT 1456 5612 1488 5644 ;
    LAYER V1 ;
      RECT 1520 152 1552 184 ;
    LAYER V1 ;
      RECT 1584 5612 1616 5644 ;
    LAYER V1 ;
      RECT 1648 152 1680 184 ;
    LAYER V1 ;
      RECT 1712 5612 1744 5644 ;
    LAYER V1 ;
      RECT 1776 152 1808 184 ;
    LAYER V1 ;
      RECT 1840 5612 1872 5644 ;
    LAYER V1 ;
      RECT 1904 152 1936 184 ;
    LAYER V1 ;
      RECT 1968 5612 2000 5644 ;
    LAYER V1 ;
      RECT 2032 152 2064 184 ;
    LAYER V1 ;
      RECT 2096 5612 2128 5644 ;
    LAYER V1 ;
      RECT 2160 152 2192 184 ;
    LAYER V1 ;
      RECT 2224 5612 2256 5644 ;
    LAYER V1 ;
      RECT 2288 152 2320 184 ;
    LAYER V1 ;
      RECT 2352 5612 2384 5644 ;
    LAYER V1 ;
      RECT 2416 152 2448 184 ;
    LAYER V1 ;
      RECT 2480 5612 2512 5644 ;
    LAYER V1 ;
      RECT 2544 152 2576 184 ;
    LAYER V1 ;
      RECT 2608 5612 2640 5644 ;
    LAYER V1 ;
      RECT 2672 152 2704 184 ;
    LAYER V1 ;
      RECT 2736 5612 2768 5644 ;
    LAYER V1 ;
      RECT 2800 152 2832 184 ;
    LAYER V1 ;
      RECT 2864 5612 2896 5644 ;
    LAYER V1 ;
      RECT 2928 152 2960 184 ;
    LAYER V1 ;
      RECT 2992 5612 3024 5644 ;
    LAYER V1 ;
      RECT 3056 152 3088 184 ;
    LAYER V1 ;
      RECT 3120 5612 3152 5644 ;
    LAYER V1 ;
      RECT 3184 152 3216 184 ;
    LAYER V1 ;
      RECT 3248 5612 3280 5644 ;
    LAYER V1 ;
      RECT 3312 152 3344 184 ;
    LAYER V1 ;
      RECT 3376 5612 3408 5644 ;
    LAYER V1 ;
      RECT 3440 152 3472 184 ;
    LAYER V1 ;
      RECT 3504 5612 3536 5644 ;
    LAYER V1 ;
      RECT 3568 152 3600 184 ;
    LAYER V1 ;
      RECT 3632 5612 3664 5644 ;
    LAYER V1 ;
      RECT 3696 152 3728 184 ;
    LAYER V1 ;
      RECT 3760 5612 3792 5644 ;
    LAYER V1 ;
      RECT 3824 152 3856 184 ;
    LAYER V1 ;
      RECT 3888 5612 3920 5644 ;
    LAYER V1 ;
      RECT 3952 152 3984 184 ;
    LAYER V1 ;
      RECT 4016 5612 4048 5644 ;
    LAYER V1 ;
      RECT 4080 152 4112 184 ;
    LAYER V1 ;
      RECT 4144 5612 4176 5644 ;
    LAYER V1 ;
      RECT 4208 152 4240 184 ;
    LAYER V1 ;
      RECT 4272 5612 4304 5644 ;
    LAYER V1 ;
      RECT 4336 152 4368 184 ;
    LAYER V1 ;
      RECT 4400 5612 4432 5644 ;
    LAYER V1 ;
      RECT 4464 152 4496 184 ;
    LAYER V1 ;
      RECT 4528 5612 4560 5644 ;
    LAYER V1 ;
      RECT 4592 152 4624 184 ;
    LAYER V1 ;
      RECT 4656 5612 4688 5644 ;
    LAYER V1 ;
      RECT 4720 152 4752 184 ;
    LAYER V1 ;
      RECT 4784 5612 4816 5644 ;
    LAYER V1 ;
      RECT 4848 152 4880 184 ;
    LAYER V1 ;
      RECT 4912 5612 4944 5644 ;
    LAYER V1 ;
      RECT 4976 152 5008 184 ;
    LAYER V1 ;
      RECT 5040 5612 5072 5644 ;
    LAYER V1 ;
      RECT 5104 152 5136 184 ;
    LAYER V1 ;
      RECT 5168 5612 5200 5644 ;
    LAYER V1 ;
      RECT 5232 152 5264 184 ;
    LAYER V1 ;
      RECT 5296 5612 5328 5644 ;
    LAYER V1 ;
      RECT 5360 152 5392 184 ;
    LAYER V1 ;
      RECT 5424 5612 5456 5644 ;
    LAYER V1 ;
      RECT 5488 152 5520 184 ;
    LAYER V1 ;
      RECT 5552 5612 5584 5644 ;
    LAYER V1 ;
      RECT 5616 152 5648 184 ;
    LAYER V1 ;
      RECT 5680 5612 5712 5644 ;
    LAYER V1 ;
      RECT 5744 152 5776 184 ;
    LAYER V1 ;
      RECT 5744 280 5776 312 ;
    LAYER V1 ;
      RECT 5744 408 5776 440 ;
    LAYER V1 ;
      RECT 5744 536 5776 568 ;
    LAYER V1 ;
      RECT 5744 664 5776 696 ;
    LAYER V1 ;
      RECT 5744 792 5776 824 ;
    LAYER V1 ;
      RECT 5744 920 5776 952 ;
    LAYER V1 ;
      RECT 5744 1048 5776 1080 ;
    LAYER V1 ;
      RECT 5744 1176 5776 1208 ;
    LAYER V1 ;
      RECT 5744 1304 5776 1336 ;
    LAYER V1 ;
      RECT 5744 1432 5776 1464 ;
    LAYER V1 ;
      RECT 5744 1560 5776 1592 ;
    LAYER V1 ;
      RECT 5744 1688 5776 1720 ;
    LAYER V1 ;
      RECT 5744 1816 5776 1848 ;
    LAYER V1 ;
      RECT 5744 1944 5776 1976 ;
    LAYER V1 ;
      RECT 5744 2072 5776 2104 ;
    LAYER V1 ;
      RECT 5744 2200 5776 2232 ;
    LAYER V1 ;
      RECT 5744 2328 5776 2360 ;
    LAYER V1 ;
      RECT 5744 2456 5776 2488 ;
    LAYER V1 ;
      RECT 5744 2584 5776 2616 ;
    LAYER V1 ;
      RECT 5744 2712 5776 2744 ;
    LAYER V1 ;
      RECT 5744 2840 5776 2872 ;
    LAYER V1 ;
      RECT 5744 2968 5776 3000 ;
    LAYER V1 ;
      RECT 5744 3096 5776 3128 ;
    LAYER V1 ;
      RECT 5744 3224 5776 3256 ;
    LAYER V1 ;
      RECT 5744 3352 5776 3384 ;
    LAYER V1 ;
      RECT 5744 3480 5776 3512 ;
    LAYER V1 ;
      RECT 5744 3608 5776 3640 ;
    LAYER V1 ;
      RECT 5744 3736 5776 3768 ;
    LAYER V1 ;
      RECT 5744 3864 5776 3896 ;
    LAYER V1 ;
      RECT 5744 3992 5776 4024 ;
    LAYER V1 ;
      RECT 5744 4120 5776 4152 ;
    LAYER V1 ;
      RECT 5744 4248 5776 4280 ;
    LAYER V1 ;
      RECT 5744 4376 5776 4408 ;
    LAYER V1 ;
      RECT 5744 4504 5776 4536 ;
    LAYER V1 ;
      RECT 5744 4632 5776 4664 ;
    LAYER V1 ;
      RECT 5744 4760 5776 4792 ;
    LAYER V1 ;
      RECT 5744 4888 5776 4920 ;
    LAYER V1 ;
      RECT 5744 5016 5776 5048 ;
    LAYER V1 ;
      RECT 5744 5144 5776 5176 ;
    LAYER V1 ;
      RECT 5744 5272 5776 5304 ;
    LAYER V1 ;
      RECT 5744 5400 5776 5432 ;
    LAYER V1 ;
      RECT 5744 5528 5776 5560 ;
    LAYER M3 ;
      RECT 304 132 336 5664 ;
    LAYER M3 ;
      RECT 368 132 400 5664 ;
    LAYER M3 ;
      RECT 432 132 464 5664 ;
    LAYER M3 ;
      RECT 496 132 528 5664 ;
    LAYER M3 ;
      RECT 560 132 592 5664 ;
    LAYER M3 ;
      RECT 624 132 656 5664 ;
    LAYER M3 ;
      RECT 688 132 720 5664 ;
    LAYER M3 ;
      RECT 752 132 784 5664 ;
    LAYER M3 ;
      RECT 816 132 848 5664 ;
    LAYER M3 ;
      RECT 880 132 912 5664 ;
    LAYER M3 ;
      RECT 944 132 976 5664 ;
    LAYER M3 ;
      RECT 1008 132 1040 5664 ;
    LAYER M3 ;
      RECT 1072 132 1104 5664 ;
    LAYER M3 ;
      RECT 1136 132 1168 5664 ;
    LAYER M3 ;
      RECT 1200 132 1232 5664 ;
    LAYER M3 ;
      RECT 1264 132 1296 5664 ;
    LAYER M3 ;
      RECT 1328 132 1360 5664 ;
    LAYER M3 ;
      RECT 1392 132 1424 5664 ;
    LAYER M3 ;
      RECT 1456 132 1488 5664 ;
    LAYER M3 ;
      RECT 1520 132 1552 5664 ;
    LAYER M3 ;
      RECT 1584 132 1616 5664 ;
    LAYER M3 ;
      RECT 1648 132 1680 5664 ;
    LAYER M3 ;
      RECT 1712 132 1744 5664 ;
    LAYER M3 ;
      RECT 1776 132 1808 5664 ;
    LAYER M3 ;
      RECT 1840 132 1872 5664 ;
    LAYER M3 ;
      RECT 1904 132 1936 5664 ;
    LAYER M3 ;
      RECT 1968 132 2000 5664 ;
    LAYER M3 ;
      RECT 2032 132 2064 5664 ;
    LAYER M3 ;
      RECT 2096 132 2128 5664 ;
    LAYER M3 ;
      RECT 2160 132 2192 5664 ;
    LAYER M3 ;
      RECT 2224 132 2256 5664 ;
    LAYER M3 ;
      RECT 2288 132 2320 5664 ;
    LAYER M3 ;
      RECT 2352 132 2384 5664 ;
    LAYER M3 ;
      RECT 2416 132 2448 5664 ;
    LAYER M3 ;
      RECT 2480 132 2512 5664 ;
    LAYER M3 ;
      RECT 2544 132 2576 5664 ;
    LAYER M3 ;
      RECT 2608 132 2640 5664 ;
    LAYER M3 ;
      RECT 2672 132 2704 5664 ;
    LAYER M3 ;
      RECT 2736 132 2768 5664 ;
    LAYER M3 ;
      RECT 2800 132 2832 5664 ;
    LAYER M3 ;
      RECT 2864 132 2896 5664 ;
    LAYER M3 ;
      RECT 2928 132 2960 5664 ;
    LAYER M3 ;
      RECT 2992 132 3024 5664 ;
    LAYER M3 ;
      RECT 3056 132 3088 5664 ;
    LAYER M3 ;
      RECT 3120 132 3152 5664 ;
    LAYER M3 ;
      RECT 3184 132 3216 5664 ;
    LAYER M3 ;
      RECT 3248 132 3280 5664 ;
    LAYER M3 ;
      RECT 3312 132 3344 5664 ;
    LAYER M3 ;
      RECT 3376 132 3408 5664 ;
    LAYER M3 ;
      RECT 3440 132 3472 5664 ;
    LAYER M3 ;
      RECT 3504 132 3536 5664 ;
    LAYER M3 ;
      RECT 3568 132 3600 5664 ;
    LAYER M3 ;
      RECT 3632 132 3664 5664 ;
    LAYER M3 ;
      RECT 3696 132 3728 5664 ;
    LAYER M3 ;
      RECT 3760 132 3792 5664 ;
    LAYER M3 ;
      RECT 3824 132 3856 5664 ;
    LAYER M3 ;
      RECT 3888 132 3920 5664 ;
    LAYER M3 ;
      RECT 3952 132 3984 5664 ;
    LAYER M3 ;
      RECT 4016 132 4048 5664 ;
    LAYER M3 ;
      RECT 4080 132 4112 5664 ;
    LAYER M3 ;
      RECT 4144 132 4176 5664 ;
    LAYER M3 ;
      RECT 4208 132 4240 5664 ;
    LAYER M3 ;
      RECT 4272 132 4304 5664 ;
    LAYER M3 ;
      RECT 4336 132 4368 5664 ;
    LAYER M3 ;
      RECT 4400 132 4432 5664 ;
    LAYER M3 ;
      RECT 4464 132 4496 5664 ;
    LAYER M3 ;
      RECT 4528 132 4560 5664 ;
    LAYER M3 ;
      RECT 4592 132 4624 5664 ;
    LAYER M3 ;
      RECT 4656 132 4688 5664 ;
    LAYER M3 ;
      RECT 4720 132 4752 5664 ;
    LAYER M3 ;
      RECT 4784 132 4816 5664 ;
    LAYER M3 ;
      RECT 4848 132 4880 5664 ;
    LAYER M3 ;
      RECT 4912 132 4944 5664 ;
    LAYER M3 ;
      RECT 4976 132 5008 5664 ;
    LAYER M3 ;
      RECT 5040 132 5072 5664 ;
    LAYER M3 ;
      RECT 5104 132 5136 5664 ;
    LAYER M3 ;
      RECT 5168 132 5200 5664 ;
    LAYER M3 ;
      RECT 5232 132 5264 5664 ;
    LAYER M3 ;
      RECT 5296 132 5328 5664 ;
    LAYER M3 ;
      RECT 5360 132 5392 5664 ;
    LAYER M3 ;
      RECT 5424 132 5456 5664 ;
    LAYER M3 ;
      RECT 5488 132 5520 5664 ;
    LAYER M3 ;
      RECT 5552 132 5584 5664 ;
    LAYER M3 ;
      RECT 5616 132 5648 5664 ;
    LAYER M3 ;
      RECT 5680 132 5712 5664 ;
    LAYER M3 ;
      RECT 5740 132 5780 5664 ;
    LAYER V2 ;
      RECT 304 216 336 248 ;
    LAYER V2 ;
      RECT 304 344 336 376 ;
    LAYER V2 ;
      RECT 304 472 336 504 ;
    LAYER V2 ;
      RECT 304 600 336 632 ;
    LAYER V2 ;
      RECT 304 728 336 760 ;
    LAYER V2 ;
      RECT 304 856 336 888 ;
    LAYER V2 ;
      RECT 304 984 336 1016 ;
    LAYER V2 ;
      RECT 304 1112 336 1144 ;
    LAYER V2 ;
      RECT 304 1240 336 1272 ;
    LAYER V2 ;
      RECT 304 1368 336 1400 ;
    LAYER V2 ;
      RECT 304 1496 336 1528 ;
    LAYER V2 ;
      RECT 304 1624 336 1656 ;
    LAYER V2 ;
      RECT 304 1752 336 1784 ;
    LAYER V2 ;
      RECT 304 1880 336 1912 ;
    LAYER V2 ;
      RECT 304 2008 336 2040 ;
    LAYER V2 ;
      RECT 304 2136 336 2168 ;
    LAYER V2 ;
      RECT 304 2264 336 2296 ;
    LAYER V2 ;
      RECT 304 2392 336 2424 ;
    LAYER V2 ;
      RECT 304 2520 336 2552 ;
    LAYER V2 ;
      RECT 304 2648 336 2680 ;
    LAYER V2 ;
      RECT 304 2776 336 2808 ;
    LAYER V2 ;
      RECT 304 2904 336 2936 ;
    LAYER V2 ;
      RECT 304 3032 336 3064 ;
    LAYER V2 ;
      RECT 304 3160 336 3192 ;
    LAYER V2 ;
      RECT 304 3288 336 3320 ;
    LAYER V2 ;
      RECT 304 3416 336 3448 ;
    LAYER V2 ;
      RECT 304 3544 336 3576 ;
    LAYER V2 ;
      RECT 304 3672 336 3704 ;
    LAYER V2 ;
      RECT 304 3800 336 3832 ;
    LAYER V2 ;
      RECT 304 3928 336 3960 ;
    LAYER V2 ;
      RECT 304 4056 336 4088 ;
    LAYER V2 ;
      RECT 304 4184 336 4216 ;
    LAYER V2 ;
      RECT 304 4312 336 4344 ;
    LAYER V2 ;
      RECT 304 4440 336 4472 ;
    LAYER V2 ;
      RECT 304 4568 336 4600 ;
    LAYER V2 ;
      RECT 304 4696 336 4728 ;
    LAYER V2 ;
      RECT 304 4824 336 4856 ;
    LAYER V2 ;
      RECT 304 4952 336 4984 ;
    LAYER V2 ;
      RECT 304 5080 336 5112 ;
    LAYER V2 ;
      RECT 304 5208 336 5240 ;
    LAYER V2 ;
      RECT 304 5336 336 5368 ;
    LAYER V2 ;
      RECT 304 5464 336 5496 ;
    LAYER V2 ;
      RECT 304 5612 336 5644 ;
    LAYER V2 ;
      RECT 368 152 400 184 ;
    LAYER V2 ;
      RECT 432 5612 464 5644 ;
    LAYER V2 ;
      RECT 496 152 528 184 ;
    LAYER V2 ;
      RECT 560 5612 592 5644 ;
    LAYER V2 ;
      RECT 624 152 656 184 ;
    LAYER V2 ;
      RECT 688 5612 720 5644 ;
    LAYER V2 ;
      RECT 752 152 784 184 ;
    LAYER V2 ;
      RECT 816 5612 848 5644 ;
    LAYER V2 ;
      RECT 880 152 912 184 ;
    LAYER V2 ;
      RECT 944 5612 976 5644 ;
    LAYER V2 ;
      RECT 1008 152 1040 184 ;
    LAYER V2 ;
      RECT 1072 5612 1104 5644 ;
    LAYER V2 ;
      RECT 1136 152 1168 184 ;
    LAYER V2 ;
      RECT 1200 5612 1232 5644 ;
    LAYER V2 ;
      RECT 1264 152 1296 184 ;
    LAYER V2 ;
      RECT 1328 5612 1360 5644 ;
    LAYER V2 ;
      RECT 1392 152 1424 184 ;
    LAYER V2 ;
      RECT 1456 5612 1488 5644 ;
    LAYER V2 ;
      RECT 1520 152 1552 184 ;
    LAYER V2 ;
      RECT 1584 5612 1616 5644 ;
    LAYER V2 ;
      RECT 1648 152 1680 184 ;
    LAYER V2 ;
      RECT 1712 5612 1744 5644 ;
    LAYER V2 ;
      RECT 1776 152 1808 184 ;
    LAYER V2 ;
      RECT 1840 5612 1872 5644 ;
    LAYER V2 ;
      RECT 1904 152 1936 184 ;
    LAYER V2 ;
      RECT 1968 5612 2000 5644 ;
    LAYER V2 ;
      RECT 2032 152 2064 184 ;
    LAYER V2 ;
      RECT 2096 5612 2128 5644 ;
    LAYER V2 ;
      RECT 2160 152 2192 184 ;
    LAYER V2 ;
      RECT 2224 5612 2256 5644 ;
    LAYER V2 ;
      RECT 2288 152 2320 184 ;
    LAYER V2 ;
      RECT 2352 5612 2384 5644 ;
    LAYER V2 ;
      RECT 2416 152 2448 184 ;
    LAYER V2 ;
      RECT 2480 5612 2512 5644 ;
    LAYER V2 ;
      RECT 2544 152 2576 184 ;
    LAYER V2 ;
      RECT 2608 5612 2640 5644 ;
    LAYER V2 ;
      RECT 2672 152 2704 184 ;
    LAYER V2 ;
      RECT 2736 5612 2768 5644 ;
    LAYER V2 ;
      RECT 2800 152 2832 184 ;
    LAYER V2 ;
      RECT 2864 5612 2896 5644 ;
    LAYER V2 ;
      RECT 2928 152 2960 184 ;
    LAYER V2 ;
      RECT 2992 5612 3024 5644 ;
    LAYER V2 ;
      RECT 3056 152 3088 184 ;
    LAYER V2 ;
      RECT 3120 5612 3152 5644 ;
    LAYER V2 ;
      RECT 3184 152 3216 184 ;
    LAYER V2 ;
      RECT 3248 5612 3280 5644 ;
    LAYER V2 ;
      RECT 3312 152 3344 184 ;
    LAYER V2 ;
      RECT 3376 5612 3408 5644 ;
    LAYER V2 ;
      RECT 3440 152 3472 184 ;
    LAYER V2 ;
      RECT 3504 5612 3536 5644 ;
    LAYER V2 ;
      RECT 3568 152 3600 184 ;
    LAYER V2 ;
      RECT 3632 5612 3664 5644 ;
    LAYER V2 ;
      RECT 3696 152 3728 184 ;
    LAYER V2 ;
      RECT 3760 5612 3792 5644 ;
    LAYER V2 ;
      RECT 3824 152 3856 184 ;
    LAYER V2 ;
      RECT 3888 5612 3920 5644 ;
    LAYER V2 ;
      RECT 3952 152 3984 184 ;
    LAYER V2 ;
      RECT 4016 5612 4048 5644 ;
    LAYER V2 ;
      RECT 4080 152 4112 184 ;
    LAYER V2 ;
      RECT 4144 5612 4176 5644 ;
    LAYER V2 ;
      RECT 4208 152 4240 184 ;
    LAYER V2 ;
      RECT 4272 5612 4304 5644 ;
    LAYER V2 ;
      RECT 4336 152 4368 184 ;
    LAYER V2 ;
      RECT 4400 5612 4432 5644 ;
    LAYER V2 ;
      RECT 4464 152 4496 184 ;
    LAYER V2 ;
      RECT 4528 5612 4560 5644 ;
    LAYER V2 ;
      RECT 4592 152 4624 184 ;
    LAYER V2 ;
      RECT 4656 5612 4688 5644 ;
    LAYER V2 ;
      RECT 4720 152 4752 184 ;
    LAYER V2 ;
      RECT 4784 5612 4816 5644 ;
    LAYER V2 ;
      RECT 4848 152 4880 184 ;
    LAYER V2 ;
      RECT 4912 5612 4944 5644 ;
    LAYER V2 ;
      RECT 4976 152 5008 184 ;
    LAYER V2 ;
      RECT 5040 5612 5072 5644 ;
    LAYER V2 ;
      RECT 5104 152 5136 184 ;
    LAYER V2 ;
      RECT 5168 5612 5200 5644 ;
    LAYER V2 ;
      RECT 5232 152 5264 184 ;
    LAYER V2 ;
      RECT 5296 5612 5328 5644 ;
    LAYER V2 ;
      RECT 5360 152 5392 184 ;
    LAYER V2 ;
      RECT 5424 5612 5456 5644 ;
    LAYER V2 ;
      RECT 5488 152 5520 184 ;
    LAYER V2 ;
      RECT 5552 5612 5584 5644 ;
    LAYER V2 ;
      RECT 5616 152 5648 184 ;
    LAYER V2 ;
      RECT 5680 5612 5712 5644 ;
    LAYER V2 ;
      RECT 5744 152 5776 184 ;
    LAYER V2 ;
      RECT 5744 280 5776 312 ;
    LAYER V2 ;
      RECT 5744 408 5776 440 ;
    LAYER V2 ;
      RECT 5744 536 5776 568 ;
    LAYER V2 ;
      RECT 5744 664 5776 696 ;
    LAYER V2 ;
      RECT 5744 792 5776 824 ;
    LAYER V2 ;
      RECT 5744 920 5776 952 ;
    LAYER V2 ;
      RECT 5744 1048 5776 1080 ;
    LAYER V2 ;
      RECT 5744 1176 5776 1208 ;
    LAYER V2 ;
      RECT 5744 1304 5776 1336 ;
    LAYER V2 ;
      RECT 5744 1432 5776 1464 ;
    LAYER V2 ;
      RECT 5744 1560 5776 1592 ;
    LAYER V2 ;
      RECT 5744 1688 5776 1720 ;
    LAYER V2 ;
      RECT 5744 1816 5776 1848 ;
    LAYER V2 ;
      RECT 5744 1944 5776 1976 ;
    LAYER V2 ;
      RECT 5744 2072 5776 2104 ;
    LAYER V2 ;
      RECT 5744 2200 5776 2232 ;
    LAYER V2 ;
      RECT 5744 2328 5776 2360 ;
    LAYER V2 ;
      RECT 5744 2456 5776 2488 ;
    LAYER V2 ;
      RECT 5744 2584 5776 2616 ;
    LAYER V2 ;
      RECT 5744 2712 5776 2744 ;
    LAYER V2 ;
      RECT 5744 2840 5776 2872 ;
    LAYER V2 ;
      RECT 5744 2968 5776 3000 ;
    LAYER V2 ;
      RECT 5744 3096 5776 3128 ;
    LAYER V2 ;
      RECT 5744 3224 5776 3256 ;
    LAYER V2 ;
      RECT 5744 3352 5776 3384 ;
    LAYER V2 ;
      RECT 5744 3480 5776 3512 ;
    LAYER V2 ;
      RECT 5744 3608 5776 3640 ;
    LAYER V2 ;
      RECT 5744 3736 5776 3768 ;
    LAYER V2 ;
      RECT 5744 3864 5776 3896 ;
    LAYER V2 ;
      RECT 5744 3992 5776 4024 ;
    LAYER V2 ;
      RECT 5744 4120 5776 4152 ;
    LAYER V2 ;
      RECT 5744 4248 5776 4280 ;
    LAYER V2 ;
      RECT 5744 4376 5776 4408 ;
    LAYER V2 ;
      RECT 5744 4504 5776 4536 ;
    LAYER V2 ;
      RECT 5744 4632 5776 4664 ;
    LAYER V2 ;
      RECT 5744 4760 5776 4792 ;
    LAYER V2 ;
      RECT 5744 4888 5776 4920 ;
    LAYER V2 ;
      RECT 5744 5016 5776 5048 ;
    LAYER V2 ;
      RECT 5744 5144 5776 5176 ;
    LAYER V2 ;
      RECT 5744 5272 5776 5304 ;
    LAYER V2 ;
      RECT 5744 5400 5776 5432 ;
    LAYER V2 ;
      RECT 5744 5528 5776 5560 ;
  END
END CAP_2T_57809468
MACRO NMOS_4T_21841201_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_4T_21841201_X1_Y1 0 0 ;
  SIZE 640 BY 2352 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124 1748 356 1780 ;
    END
  END B
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124 68 356 100 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124 908 356 940 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204 152 436 184 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1644 336 1884 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1748 336 1780 ;
    LAYER V1 ;
      RECT 224 152 256 184 ;
    LAYER V1 ;
      RECT 384 152 416 184 ;
    LAYER V0 ;
      RECT 304 461 336 493 ;
    LAYER V0 ;
      RECT 304 545 336 577 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1748 336 1780 ;
    LAYER V0 ;
      RECT 224 461 256 493 ;
    LAYER V0 ;
      RECT 224 545 256 577 ;
    LAYER V0 ;
      RECT 384 461 416 493 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
  END
END NMOS_4T_21841201_X1_Y1
MACRO PMOS_S_32697230_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN PMOS_S_32697230_X1_Y1 0 0 ;
  SIZE 640 BY 2352 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124 68 356 100 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124 908 356 940 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 220 132 260 1800 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1644 336 1884 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M2 ;
      RECT 124 1748 356 1780 ;
    LAYER M2 ;
      RECT 204 152 436 184 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1748 336 1780 ;
    LAYER V1 ;
      RECT 224 152 256 184 ;
    LAYER V1 ;
      RECT 384 152 416 184 ;
    LAYER V2 ;
      RECT 224 152 256 184 ;
    LAYER V2 ;
      RECT 224 1748 256 1780 ;
    LAYER V0 ;
      RECT 304 335 336 367 ;
    LAYER V0 ;
      RECT 304 419 336 451 ;
    LAYER V0 ;
      RECT 304 503 336 535 ;
    LAYER V0 ;
      RECT 304 587 336 619 ;
    LAYER V0 ;
      RECT 304 671 336 703 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1748 336 1780 ;
    LAYER V0 ;
      RECT 224 335 256 367 ;
    LAYER V0 ;
      RECT 224 419 256 451 ;
    LAYER V0 ;
      RECT 224 503 256 535 ;
    LAYER V0 ;
      RECT 224 587 256 619 ;
    LAYER V0 ;
      RECT 224 671 256 703 ;
    LAYER V0 ;
      RECT 384 335 416 367 ;
    LAYER V0 ;
      RECT 384 419 416 451 ;
    LAYER V0 ;
      RECT 384 503 416 535 ;
    LAYER V0 ;
      RECT 384 587 416 619 ;
    LAYER V0 ;
      RECT 384 671 416 703 ;
  END
END PMOS_S_32697230_X1_Y1
