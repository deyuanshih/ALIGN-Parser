MACRO CCP_NMOS_23282412_X2_Y2
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CCP_NMOS_23282412_X2_Y2 0 0 ;
  SIZE 1120 BY 3528 ;
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 300 48 340 2136 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 380 132 420 2220 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 460 216 500 2976 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1224 336 1968 ;
    LAYER M1 ;
      RECT 304 2064 336 2304 ;
    LAYER M1 ;
      RECT 304 2820 336 3060 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 224 1224 256 1968 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 384 1224 416 1968 ;
    LAYER M1 ;
      RECT 464 48 496 792 ;
    LAYER M1 ;
      RECT 464 888 496 1128 ;
    LAYER M1 ;
      RECT 464 1224 496 1968 ;
    LAYER M1 ;
      RECT 464 2064 496 2304 ;
    LAYER M1 ;
      RECT 464 2820 496 3060 ;
    LAYER M1 ;
      RECT 544 48 576 792 ;
    LAYER M1 ;
      RECT 544 1224 576 1968 ;
    LAYER M1 ;
      RECT 624 48 656 792 ;
    LAYER M1 ;
      RECT 624 888 656 1128 ;
    LAYER M1 ;
      RECT 624 1224 656 1968 ;
    LAYER M1 ;
      RECT 624 2064 656 2304 ;
    LAYER M1 ;
      RECT 624 2820 656 3060 ;
    LAYER M1 ;
      RECT 704 48 736 792 ;
    LAYER M1 ;
      RECT 704 1224 736 1968 ;
    LAYER M1 ;
      RECT 784 48 816 792 ;
    LAYER M1 ;
      RECT 784 888 816 1128 ;
    LAYER M1 ;
      RECT 784 1224 816 1968 ;
    LAYER M1 ;
      RECT 784 2064 816 2304 ;
    LAYER M1 ;
      RECT 784 2820 816 3060 ;
    LAYER M1 ;
      RECT 864 48 896 792 ;
    LAYER M1 ;
      RECT 864 1224 896 1968 ;
    LAYER M2 ;
      RECT 284 908 676 940 ;
    LAYER M2 ;
      RECT 284 68 836 100 ;
    LAYER M2 ;
      RECT 284 992 836 1024 ;
    LAYER M2 ;
      RECT 364 152 676 184 ;
    LAYER M2 ;
      RECT 204 236 916 268 ;
    LAYER M2 ;
      RECT 284 2084 836 2116 ;
    LAYER M2 ;
      RECT 284 1244 676 1276 ;
    LAYER M2 ;
      RECT 364 2168 676 2200 ;
    LAYER M2 ;
      RECT 284 1328 836 1360 ;
    LAYER M2 ;
      RECT 284 2924 836 2956 ;
    LAYER M2 ;
      RECT 204 1412 916 1444 ;
    LAYER V1 ;
      RECT 624 152 656 184 ;
    LAYER V1 ;
      RECT 624 908 656 940 ;
    LAYER V1 ;
      RECT 624 1244 656 1276 ;
    LAYER V1 ;
      RECT 624 2168 656 2200 ;
    LAYER V1 ;
      RECT 624 2924 656 2956 ;
    LAYER V1 ;
      RECT 464 152 496 184 ;
    LAYER V1 ;
      RECT 464 908 496 940 ;
    LAYER V1 ;
      RECT 464 1244 496 1276 ;
    LAYER V1 ;
      RECT 464 2168 496 2200 ;
    LAYER V1 ;
      RECT 464 2924 496 2956 ;
    LAYER V1 ;
      RECT 784 68 816 100 ;
    LAYER V1 ;
      RECT 784 992 816 1024 ;
    LAYER V1 ;
      RECT 784 1328 816 1360 ;
    LAYER V1 ;
      RECT 784 2084 816 2116 ;
    LAYER V1 ;
      RECT 784 2924 816 2956 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 992 336 1024 ;
    LAYER V1 ;
      RECT 304 1328 336 1360 ;
    LAYER V1 ;
      RECT 304 2084 336 2116 ;
    LAYER V1 ;
      RECT 304 2924 336 2956 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 224 1412 256 1444 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 384 1412 416 1444 ;
    LAYER V1 ;
      RECT 544 236 576 268 ;
    LAYER V1 ;
      RECT 544 1412 576 1444 ;
    LAYER V1 ;
      RECT 704 236 736 268 ;
    LAYER V1 ;
      RECT 704 1412 736 1444 ;
    LAYER V1 ;
      RECT 864 236 896 268 ;
    LAYER V1 ;
      RECT 864 1412 896 1444 ;
    LAYER V2 ;
      RECT 304 68 336 100 ;
    LAYER V2 ;
      RECT 304 908 336 940 ;
    LAYER V2 ;
      RECT 304 1244 336 1276 ;
    LAYER V2 ;
      RECT 304 2084 336 2116 ;
    LAYER V2 ;
      RECT 384 152 416 184 ;
    LAYER V2 ;
      RECT 384 992 416 1024 ;
    LAYER V2 ;
      RECT 384 1328 416 1360 ;
    LAYER V2 ;
      RECT 384 2168 416 2200 ;
    LAYER V2 ;
      RECT 464 236 496 268 ;
    LAYER V2 ;
      RECT 464 1412 496 1444 ;
    LAYER V2 ;
      RECT 464 2924 496 2956 ;
    LAYER V0 ;
      RECT 304 545 336 577 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1721 336 1753 ;
    LAYER V0 ;
      RECT 304 2084 336 2116 ;
    LAYER V0 ;
      RECT 304 2924 336 2956 ;
    LAYER V0 ;
      RECT 304 2924 336 2956 ;
    LAYER V0 ;
      RECT 224 545 256 577 ;
    LAYER V0 ;
      RECT 224 1721 256 1753 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 384 1721 416 1753 ;
    LAYER V0 ;
      RECT 384 1721 416 1753 ;
    LAYER V0 ;
      RECT 464 545 496 577 ;
    LAYER V0 ;
      RECT 464 908 496 940 ;
    LAYER V0 ;
      RECT 464 1721 496 1753 ;
    LAYER V0 ;
      RECT 464 2084 496 2116 ;
    LAYER V0 ;
      RECT 464 2924 496 2956 ;
    LAYER V0 ;
      RECT 464 2924 496 2956 ;
    LAYER V0 ;
      RECT 544 545 576 577 ;
    LAYER V0 ;
      RECT 544 545 576 577 ;
    LAYER V0 ;
      RECT 544 1721 576 1753 ;
    LAYER V0 ;
      RECT 544 1721 576 1753 ;
    LAYER V0 ;
      RECT 624 545 656 577 ;
    LAYER V0 ;
      RECT 624 908 656 940 ;
    LAYER V0 ;
      RECT 624 1721 656 1753 ;
    LAYER V0 ;
      RECT 624 2084 656 2116 ;
    LAYER V0 ;
      RECT 624 2924 656 2956 ;
    LAYER V0 ;
      RECT 624 2924 656 2956 ;
    LAYER V0 ;
      RECT 704 545 736 577 ;
    LAYER V0 ;
      RECT 704 545 736 577 ;
    LAYER V0 ;
      RECT 704 1721 736 1753 ;
    LAYER V0 ;
      RECT 704 1721 736 1753 ;
    LAYER V0 ;
      RECT 784 545 816 577 ;
    LAYER V0 ;
      RECT 784 908 816 940 ;
    LAYER V0 ;
      RECT 784 1721 816 1753 ;
    LAYER V0 ;
      RECT 784 2084 816 2116 ;
    LAYER V0 ;
      RECT 784 2924 816 2956 ;
    LAYER V0 ;
      RECT 784 2924 816 2956 ;
    LAYER V0 ;
      RECT 864 545 896 577 ;
    LAYER V0 ;
      RECT 864 1721 896 1753 ;
  END
END CCP_NMOS_23282412_X2_Y2
