MACRO CMC_S_PMOS_70942995
  ORIGIN 0 0 ;
  FOREIGN CMC_S_PMOS_70942995 0 0 ;
  SIZE 1.28 BY 2.352 ;
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.284 0.068 0.516 0.1 ;
    END
  END DA
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.284 0.908 0.516 0.94 ;
      LAYER M2 ;
        RECT 0.764 0.908 0.996 0.94 ;
      LAYER M2 ;
        RECT 0.48 0.908 0.8 0.94 ;
    END
  END G
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 0.38 0.132 0.42 1.8 ;
    END
  END SA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.764 0.068 0.996 0.1 ;
    END
  END DB
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 0.86 0.132 0.9 1.8 ;
    END
  END SB
  OBS 
  LAYER M1 ;
        RECT 0.304 0.048 0.336 0.792 ;
  LAYER M1 ;
        RECT 0.304 0.888 0.336 1.128 ;
  LAYER M1 ;
        RECT 0.304 1.644 0.336 1.884 ;
  LAYER M1 ;
        RECT 0.384 0.048 0.416 0.792 ;
  LAYER M1 ;
        RECT 0.224 0.048 0.256 0.792 ;
  LAYER M2 ;
        RECT 0.284 1.748 0.516 1.78 ;
  LAYER M2 ;
        RECT 0.204 0.152 0.436 0.184 ;
  LAYER M2 ;
        RECT 0.284 0.068 0.516 0.1 ;
  LAYER M2 ;
        RECT 0.284 0.908 0.516 0.94 ;
  LAYER M3 ;
        RECT 0.38 0.132 0.42 1.8 ;
  LAYER M1 ;
        RECT 0.944 0.048 0.976 0.792 ;
  LAYER M1 ;
        RECT 0.944 0.888 0.976 1.128 ;
  LAYER M1 ;
        RECT 0.944 1.644 0.976 1.884 ;
  LAYER M1 ;
        RECT 0.864 0.048 0.896 0.792 ;
  LAYER M1 ;
        RECT 1.024 0.048 1.056 0.792 ;
  LAYER M2 ;
        RECT 0.764 1.748 0.996 1.78 ;
  LAYER M2 ;
        RECT 0.844 0.152 1.076 0.184 ;
  LAYER M2 ;
        RECT 0.764 0.068 0.996 0.1 ;
  LAYER M2 ;
        RECT 0.764 0.908 0.996 0.94 ;
  LAYER M3 ;
        RECT 0.86 0.132 0.9 1.8 ;
  END 
END CMC_S_PMOS_70942995
