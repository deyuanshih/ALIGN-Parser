MACRO CAP_2T_8193393
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CAP_2T_8193393 0 0 ;
  SIZE 4480 BY 4116 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44 3932 4436 3964 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44 152 4436 184 ;
    END
  END PLUS
  OBS
    LAYER M1 ;
      RECT 304 132 336 3984 ;
    LAYER M1 ;
      RECT 368 132 400 3984 ;
    LAYER M1 ;
      RECT 432 132 464 3984 ;
    LAYER M1 ;
      RECT 496 132 528 3984 ;
    LAYER M1 ;
      RECT 560 132 592 3984 ;
    LAYER M1 ;
      RECT 624 132 656 3984 ;
    LAYER M1 ;
      RECT 688 132 720 3984 ;
    LAYER M1 ;
      RECT 752 132 784 3984 ;
    LAYER M1 ;
      RECT 816 132 848 3984 ;
    LAYER M1 ;
      RECT 880 132 912 3984 ;
    LAYER M1 ;
      RECT 944 132 976 3984 ;
    LAYER M1 ;
      RECT 1008 132 1040 3984 ;
    LAYER M1 ;
      RECT 1072 132 1104 3984 ;
    LAYER M1 ;
      RECT 1136 132 1168 3984 ;
    LAYER M1 ;
      RECT 1200 132 1232 3984 ;
    LAYER M1 ;
      RECT 1264 132 1296 3984 ;
    LAYER M1 ;
      RECT 1328 132 1360 3984 ;
    LAYER M1 ;
      RECT 1392 132 1424 3984 ;
    LAYER M1 ;
      RECT 1456 132 1488 3984 ;
    LAYER M1 ;
      RECT 1520 132 1552 3984 ;
    LAYER M1 ;
      RECT 1584 132 1616 3984 ;
    LAYER M1 ;
      RECT 1648 132 1680 3984 ;
    LAYER M1 ;
      RECT 1712 132 1744 3984 ;
    LAYER M1 ;
      RECT 1776 132 1808 3984 ;
    LAYER M1 ;
      RECT 1840 132 1872 3984 ;
    LAYER M1 ;
      RECT 1904 132 1936 3984 ;
    LAYER M1 ;
      RECT 1968 132 2000 3984 ;
    LAYER M1 ;
      RECT 2032 132 2064 3984 ;
    LAYER M1 ;
      RECT 2096 132 2128 3984 ;
    LAYER M1 ;
      RECT 2160 132 2192 3984 ;
    LAYER M1 ;
      RECT 2224 132 2256 3984 ;
    LAYER M1 ;
      RECT 2288 132 2320 3984 ;
    LAYER M1 ;
      RECT 2352 132 2384 3984 ;
    LAYER M1 ;
      RECT 2416 132 2448 3984 ;
    LAYER M1 ;
      RECT 2480 132 2512 3984 ;
    LAYER M1 ;
      RECT 2544 132 2576 3984 ;
    LAYER M1 ;
      RECT 2608 132 2640 3984 ;
    LAYER M1 ;
      RECT 2672 132 2704 3984 ;
    LAYER M1 ;
      RECT 2736 132 2768 3984 ;
    LAYER M1 ;
      RECT 2800 132 2832 3984 ;
    LAYER M1 ;
      RECT 2864 132 2896 3984 ;
    LAYER M1 ;
      RECT 2928 132 2960 3984 ;
    LAYER M1 ;
      RECT 2992 132 3024 3984 ;
    LAYER M1 ;
      RECT 3056 132 3088 3984 ;
    LAYER M1 ;
      RECT 3120 132 3152 3984 ;
    LAYER M1 ;
      RECT 3184 132 3216 3984 ;
    LAYER M1 ;
      RECT 3248 132 3280 3984 ;
    LAYER M1 ;
      RECT 3312 132 3344 3984 ;
    LAYER M1 ;
      RECT 3376 132 3408 3984 ;
    LAYER M1 ;
      RECT 3440 132 3472 3984 ;
    LAYER M1 ;
      RECT 3504 132 3536 3984 ;
    LAYER M1 ;
      RECT 3568 132 3600 3984 ;
    LAYER M1 ;
      RECT 3632 132 3664 3984 ;
    LAYER M1 ;
      RECT 3696 132 3728 3984 ;
    LAYER M1 ;
      RECT 3760 132 3792 3984 ;
    LAYER M1 ;
      RECT 3824 132 3856 3984 ;
    LAYER M1 ;
      RECT 3888 132 3920 3984 ;
    LAYER M1 ;
      RECT 3952 132 3984 3984 ;
    LAYER M1 ;
      RECT 4016 132 4048 3984 ;
    LAYER M1 ;
      RECT 4144 132 4176 3984 ;
    LAYER M2 ;
      RECT 284 216 4196 248 ;
    LAYER M2 ;
      RECT 284 280 4196 312 ;
    LAYER M2 ;
      RECT 284 344 4196 376 ;
    LAYER M2 ;
      RECT 284 408 4196 440 ;
    LAYER M2 ;
      RECT 284 472 4196 504 ;
    LAYER M2 ;
      RECT 284 536 4196 568 ;
    LAYER M2 ;
      RECT 284 600 4196 632 ;
    LAYER M2 ;
      RECT 284 664 4196 696 ;
    LAYER M2 ;
      RECT 284 728 4196 760 ;
    LAYER M2 ;
      RECT 284 792 4196 824 ;
    LAYER M2 ;
      RECT 284 856 4196 888 ;
    LAYER M2 ;
      RECT 284 920 4196 952 ;
    LAYER M2 ;
      RECT 284 984 4196 1016 ;
    LAYER M2 ;
      RECT 284 1048 4196 1080 ;
    LAYER M2 ;
      RECT 284 1112 4196 1144 ;
    LAYER M2 ;
      RECT 284 1176 4196 1208 ;
    LAYER M2 ;
      RECT 284 1240 4196 1272 ;
    LAYER M2 ;
      RECT 284 1304 4196 1336 ;
    LAYER M2 ;
      RECT 284 1368 4196 1400 ;
    LAYER M2 ;
      RECT 284 1432 4196 1464 ;
    LAYER M2 ;
      RECT 284 1496 4196 1528 ;
    LAYER M2 ;
      RECT 284 1560 4196 1592 ;
    LAYER M2 ;
      RECT 284 1624 4196 1656 ;
    LAYER M2 ;
      RECT 284 1688 4196 1720 ;
    LAYER M2 ;
      RECT 284 1752 4196 1784 ;
    LAYER M2 ;
      RECT 284 1816 4196 1848 ;
    LAYER M2 ;
      RECT 284 1880 4196 1912 ;
    LAYER M2 ;
      RECT 284 1944 4196 1976 ;
    LAYER M2 ;
      RECT 284 2008 4196 2040 ;
    LAYER M2 ;
      RECT 284 2072 4196 2104 ;
    LAYER M2 ;
      RECT 284 2136 4196 2168 ;
    LAYER M2 ;
      RECT 284 2200 4196 2232 ;
    LAYER M2 ;
      RECT 284 2264 4196 2296 ;
    LAYER M2 ;
      RECT 284 2328 4196 2360 ;
    LAYER M2 ;
      RECT 284 2392 4196 2424 ;
    LAYER M2 ;
      RECT 284 2456 4196 2488 ;
    LAYER M2 ;
      RECT 284 2520 4196 2552 ;
    LAYER M2 ;
      RECT 284 2584 4196 2616 ;
    LAYER M2 ;
      RECT 284 2648 4196 2680 ;
    LAYER M2 ;
      RECT 284 2712 4196 2744 ;
    LAYER M2 ;
      RECT 284 2776 4196 2808 ;
    LAYER M2 ;
      RECT 284 2840 4196 2872 ;
    LAYER M2 ;
      RECT 284 2904 4196 2936 ;
    LAYER M2 ;
      RECT 284 2968 4196 3000 ;
    LAYER M2 ;
      RECT 284 3032 4196 3064 ;
    LAYER M2 ;
      RECT 284 3096 4196 3128 ;
    LAYER M2 ;
      RECT 284 3160 4196 3192 ;
    LAYER M2 ;
      RECT 284 3224 4196 3256 ;
    LAYER M2 ;
      RECT 284 3288 4196 3320 ;
    LAYER M2 ;
      RECT 284 3352 4196 3384 ;
    LAYER M2 ;
      RECT 284 3416 4196 3448 ;
    LAYER M2 ;
      RECT 284 3480 4196 3512 ;
    LAYER M2 ;
      RECT 284 3544 4196 3576 ;
    LAYER M2 ;
      RECT 284 3608 4196 3640 ;
    LAYER M2 ;
      RECT 284 3672 4196 3704 ;
    LAYER M2 ;
      RECT 284 3736 4196 3768 ;
    LAYER M2 ;
      RECT 284 3800 4196 3832 ;
    LAYER M2 ;
      RECT 284 3864 4196 3896 ;
    LAYER V1 ;
      RECT 304 216 336 248 ;
    LAYER V1 ;
      RECT 304 344 336 376 ;
    LAYER V1 ;
      RECT 304 472 336 504 ;
    LAYER V1 ;
      RECT 304 600 336 632 ;
    LAYER V1 ;
      RECT 304 728 336 760 ;
    LAYER V1 ;
      RECT 304 856 336 888 ;
    LAYER V1 ;
      RECT 304 984 336 1016 ;
    LAYER V1 ;
      RECT 304 1112 336 1144 ;
    LAYER V1 ;
      RECT 304 1240 336 1272 ;
    LAYER V1 ;
      RECT 304 1368 336 1400 ;
    LAYER V1 ;
      RECT 304 1496 336 1528 ;
    LAYER V1 ;
      RECT 304 1624 336 1656 ;
    LAYER V1 ;
      RECT 304 1752 336 1784 ;
    LAYER V1 ;
      RECT 304 1880 336 1912 ;
    LAYER V1 ;
      RECT 304 2008 336 2040 ;
    LAYER V1 ;
      RECT 304 2136 336 2168 ;
    LAYER V1 ;
      RECT 304 2264 336 2296 ;
    LAYER V1 ;
      RECT 304 2392 336 2424 ;
    LAYER V1 ;
      RECT 304 2520 336 2552 ;
    LAYER V1 ;
      RECT 304 2648 336 2680 ;
    LAYER V1 ;
      RECT 304 2776 336 2808 ;
    LAYER V1 ;
      RECT 304 2904 336 2936 ;
    LAYER V1 ;
      RECT 304 3032 336 3064 ;
    LAYER V1 ;
      RECT 304 3160 336 3192 ;
    LAYER V1 ;
      RECT 304 3288 336 3320 ;
    LAYER V1 ;
      RECT 304 3416 336 3448 ;
    LAYER V1 ;
      RECT 304 3544 336 3576 ;
    LAYER V1 ;
      RECT 304 3672 336 3704 ;
    LAYER V1 ;
      RECT 304 3800 336 3832 ;
    LAYER V1 ;
      RECT 304 3932 336 3964 ;
    LAYER V1 ;
      RECT 368 152 400 184 ;
    LAYER V1 ;
      RECT 432 3932 464 3964 ;
    LAYER V1 ;
      RECT 496 152 528 184 ;
    LAYER V1 ;
      RECT 560 3932 592 3964 ;
    LAYER V1 ;
      RECT 624 152 656 184 ;
    LAYER V1 ;
      RECT 688 3932 720 3964 ;
    LAYER V1 ;
      RECT 752 152 784 184 ;
    LAYER V1 ;
      RECT 816 3932 848 3964 ;
    LAYER V1 ;
      RECT 880 152 912 184 ;
    LAYER V1 ;
      RECT 944 3932 976 3964 ;
    LAYER V1 ;
      RECT 1008 152 1040 184 ;
    LAYER V1 ;
      RECT 1072 3932 1104 3964 ;
    LAYER V1 ;
      RECT 1136 152 1168 184 ;
    LAYER V1 ;
      RECT 1200 3932 1232 3964 ;
    LAYER V1 ;
      RECT 1264 152 1296 184 ;
    LAYER V1 ;
      RECT 1328 3932 1360 3964 ;
    LAYER V1 ;
      RECT 1392 152 1424 184 ;
    LAYER V1 ;
      RECT 1456 3932 1488 3964 ;
    LAYER V1 ;
      RECT 1520 152 1552 184 ;
    LAYER V1 ;
      RECT 1584 3932 1616 3964 ;
    LAYER V1 ;
      RECT 1648 152 1680 184 ;
    LAYER V1 ;
      RECT 1712 3932 1744 3964 ;
    LAYER V1 ;
      RECT 1776 152 1808 184 ;
    LAYER V1 ;
      RECT 1840 3932 1872 3964 ;
    LAYER V1 ;
      RECT 1904 152 1936 184 ;
    LAYER V1 ;
      RECT 1968 3932 2000 3964 ;
    LAYER V1 ;
      RECT 2032 152 2064 184 ;
    LAYER V1 ;
      RECT 2096 3932 2128 3964 ;
    LAYER V1 ;
      RECT 2160 152 2192 184 ;
    LAYER V1 ;
      RECT 2224 3932 2256 3964 ;
    LAYER V1 ;
      RECT 2288 152 2320 184 ;
    LAYER V1 ;
      RECT 2352 3932 2384 3964 ;
    LAYER V1 ;
      RECT 2416 152 2448 184 ;
    LAYER V1 ;
      RECT 2480 3932 2512 3964 ;
    LAYER V1 ;
      RECT 2544 152 2576 184 ;
    LAYER V1 ;
      RECT 2608 3932 2640 3964 ;
    LAYER V1 ;
      RECT 2672 152 2704 184 ;
    LAYER V1 ;
      RECT 2736 3932 2768 3964 ;
    LAYER V1 ;
      RECT 2800 152 2832 184 ;
    LAYER V1 ;
      RECT 2864 3932 2896 3964 ;
    LAYER V1 ;
      RECT 2928 152 2960 184 ;
    LAYER V1 ;
      RECT 2992 3932 3024 3964 ;
    LAYER V1 ;
      RECT 3056 152 3088 184 ;
    LAYER V1 ;
      RECT 3120 3932 3152 3964 ;
    LAYER V1 ;
      RECT 3184 152 3216 184 ;
    LAYER V1 ;
      RECT 3248 3932 3280 3964 ;
    LAYER V1 ;
      RECT 3312 152 3344 184 ;
    LAYER V1 ;
      RECT 3376 3932 3408 3964 ;
    LAYER V1 ;
      RECT 3440 152 3472 184 ;
    LAYER V1 ;
      RECT 3504 3932 3536 3964 ;
    LAYER V1 ;
      RECT 3568 152 3600 184 ;
    LAYER V1 ;
      RECT 3632 3932 3664 3964 ;
    LAYER V1 ;
      RECT 3696 152 3728 184 ;
    LAYER V1 ;
      RECT 3760 3932 3792 3964 ;
    LAYER V1 ;
      RECT 3824 152 3856 184 ;
    LAYER V1 ;
      RECT 3888 3932 3920 3964 ;
    LAYER V1 ;
      RECT 3952 152 3984 184 ;
    LAYER V1 ;
      RECT 4016 3932 4048 3964 ;
    LAYER V1 ;
      RECT 4144 152 4176 184 ;
    LAYER V1 ;
      RECT 4144 280 4176 312 ;
    LAYER V1 ;
      RECT 4144 408 4176 440 ;
    LAYER V1 ;
      RECT 4144 536 4176 568 ;
    LAYER V1 ;
      RECT 4144 664 4176 696 ;
    LAYER V1 ;
      RECT 4144 792 4176 824 ;
    LAYER V1 ;
      RECT 4144 920 4176 952 ;
    LAYER V1 ;
      RECT 4144 1048 4176 1080 ;
    LAYER V1 ;
      RECT 4144 1176 4176 1208 ;
    LAYER V1 ;
      RECT 4144 1304 4176 1336 ;
    LAYER V1 ;
      RECT 4144 1432 4176 1464 ;
    LAYER V1 ;
      RECT 4144 1560 4176 1592 ;
    LAYER V1 ;
      RECT 4144 1688 4176 1720 ;
    LAYER V1 ;
      RECT 4144 1816 4176 1848 ;
    LAYER V1 ;
      RECT 4144 1944 4176 1976 ;
    LAYER V1 ;
      RECT 4144 2072 4176 2104 ;
    LAYER V1 ;
      RECT 4144 2200 4176 2232 ;
    LAYER V1 ;
      RECT 4144 2328 4176 2360 ;
    LAYER V1 ;
      RECT 4144 2456 4176 2488 ;
    LAYER V1 ;
      RECT 4144 2584 4176 2616 ;
    LAYER V1 ;
      RECT 4144 2712 4176 2744 ;
    LAYER V1 ;
      RECT 4144 2840 4176 2872 ;
    LAYER V1 ;
      RECT 4144 2968 4176 3000 ;
    LAYER V1 ;
      RECT 4144 3096 4176 3128 ;
    LAYER V1 ;
      RECT 4144 3224 4176 3256 ;
    LAYER V1 ;
      RECT 4144 3352 4176 3384 ;
    LAYER V1 ;
      RECT 4144 3480 4176 3512 ;
    LAYER V1 ;
      RECT 4144 3608 4176 3640 ;
    LAYER V1 ;
      RECT 4144 3736 4176 3768 ;
    LAYER V1 ;
      RECT 4144 3864 4176 3896 ;
    LAYER M3 ;
      RECT 304 132 336 3984 ;
    LAYER M3 ;
      RECT 368 132 400 3984 ;
    LAYER M3 ;
      RECT 432 132 464 3984 ;
    LAYER M3 ;
      RECT 496 132 528 3984 ;
    LAYER M3 ;
      RECT 560 132 592 3984 ;
    LAYER M3 ;
      RECT 624 132 656 3984 ;
    LAYER M3 ;
      RECT 688 132 720 3984 ;
    LAYER M3 ;
      RECT 752 132 784 3984 ;
    LAYER M3 ;
      RECT 816 132 848 3984 ;
    LAYER M3 ;
      RECT 880 132 912 3984 ;
    LAYER M3 ;
      RECT 944 132 976 3984 ;
    LAYER M3 ;
      RECT 1008 132 1040 3984 ;
    LAYER M3 ;
      RECT 1072 132 1104 3984 ;
    LAYER M3 ;
      RECT 1136 132 1168 3984 ;
    LAYER M3 ;
      RECT 1200 132 1232 3984 ;
    LAYER M3 ;
      RECT 1264 132 1296 3984 ;
    LAYER M3 ;
      RECT 1328 132 1360 3984 ;
    LAYER M3 ;
      RECT 1392 132 1424 3984 ;
    LAYER M3 ;
      RECT 1456 132 1488 3984 ;
    LAYER M3 ;
      RECT 1520 132 1552 3984 ;
    LAYER M3 ;
      RECT 1584 132 1616 3984 ;
    LAYER M3 ;
      RECT 1648 132 1680 3984 ;
    LAYER M3 ;
      RECT 1712 132 1744 3984 ;
    LAYER M3 ;
      RECT 1776 132 1808 3984 ;
    LAYER M3 ;
      RECT 1840 132 1872 3984 ;
    LAYER M3 ;
      RECT 1904 132 1936 3984 ;
    LAYER M3 ;
      RECT 1968 132 2000 3984 ;
    LAYER M3 ;
      RECT 2032 132 2064 3984 ;
    LAYER M3 ;
      RECT 2096 132 2128 3984 ;
    LAYER M3 ;
      RECT 2160 132 2192 3984 ;
    LAYER M3 ;
      RECT 2224 132 2256 3984 ;
    LAYER M3 ;
      RECT 2288 132 2320 3984 ;
    LAYER M3 ;
      RECT 2352 132 2384 3984 ;
    LAYER M3 ;
      RECT 2416 132 2448 3984 ;
    LAYER M3 ;
      RECT 2480 132 2512 3984 ;
    LAYER M3 ;
      RECT 2544 132 2576 3984 ;
    LAYER M3 ;
      RECT 2608 132 2640 3984 ;
    LAYER M3 ;
      RECT 2672 132 2704 3984 ;
    LAYER M3 ;
      RECT 2736 132 2768 3984 ;
    LAYER M3 ;
      RECT 2800 132 2832 3984 ;
    LAYER M3 ;
      RECT 2864 132 2896 3984 ;
    LAYER M3 ;
      RECT 2928 132 2960 3984 ;
    LAYER M3 ;
      RECT 2992 132 3024 3984 ;
    LAYER M3 ;
      RECT 3056 132 3088 3984 ;
    LAYER M3 ;
      RECT 3120 132 3152 3984 ;
    LAYER M3 ;
      RECT 3184 132 3216 3984 ;
    LAYER M3 ;
      RECT 3248 132 3280 3984 ;
    LAYER M3 ;
      RECT 3312 132 3344 3984 ;
    LAYER M3 ;
      RECT 3376 132 3408 3984 ;
    LAYER M3 ;
      RECT 3440 132 3472 3984 ;
    LAYER M3 ;
      RECT 3504 132 3536 3984 ;
    LAYER M3 ;
      RECT 3568 132 3600 3984 ;
    LAYER M3 ;
      RECT 3632 132 3664 3984 ;
    LAYER M3 ;
      RECT 3696 132 3728 3984 ;
    LAYER M3 ;
      RECT 3760 132 3792 3984 ;
    LAYER M3 ;
      RECT 3824 132 3856 3984 ;
    LAYER M3 ;
      RECT 3888 132 3920 3984 ;
    LAYER M3 ;
      RECT 3952 132 3984 3984 ;
    LAYER M3 ;
      RECT 4016 132 4048 3984 ;
    LAYER M3 ;
      RECT 4140 132 4180 3984 ;
    LAYER V2 ;
      RECT 304 216 336 248 ;
    LAYER V2 ;
      RECT 304 344 336 376 ;
    LAYER V2 ;
      RECT 304 472 336 504 ;
    LAYER V2 ;
      RECT 304 600 336 632 ;
    LAYER V2 ;
      RECT 304 728 336 760 ;
    LAYER V2 ;
      RECT 304 856 336 888 ;
    LAYER V2 ;
      RECT 304 984 336 1016 ;
    LAYER V2 ;
      RECT 304 1112 336 1144 ;
    LAYER V2 ;
      RECT 304 1240 336 1272 ;
    LAYER V2 ;
      RECT 304 1368 336 1400 ;
    LAYER V2 ;
      RECT 304 1496 336 1528 ;
    LAYER V2 ;
      RECT 304 1624 336 1656 ;
    LAYER V2 ;
      RECT 304 1752 336 1784 ;
    LAYER V2 ;
      RECT 304 1880 336 1912 ;
    LAYER V2 ;
      RECT 304 2008 336 2040 ;
    LAYER V2 ;
      RECT 304 2136 336 2168 ;
    LAYER V2 ;
      RECT 304 2264 336 2296 ;
    LAYER V2 ;
      RECT 304 2392 336 2424 ;
    LAYER V2 ;
      RECT 304 2520 336 2552 ;
    LAYER V2 ;
      RECT 304 2648 336 2680 ;
    LAYER V2 ;
      RECT 304 2776 336 2808 ;
    LAYER V2 ;
      RECT 304 2904 336 2936 ;
    LAYER V2 ;
      RECT 304 3032 336 3064 ;
    LAYER V2 ;
      RECT 304 3160 336 3192 ;
    LAYER V2 ;
      RECT 304 3288 336 3320 ;
    LAYER V2 ;
      RECT 304 3416 336 3448 ;
    LAYER V2 ;
      RECT 304 3544 336 3576 ;
    LAYER V2 ;
      RECT 304 3672 336 3704 ;
    LAYER V2 ;
      RECT 304 3800 336 3832 ;
    LAYER V2 ;
      RECT 304 3932 336 3964 ;
    LAYER V2 ;
      RECT 368 152 400 184 ;
    LAYER V2 ;
      RECT 432 3932 464 3964 ;
    LAYER V2 ;
      RECT 496 152 528 184 ;
    LAYER V2 ;
      RECT 560 3932 592 3964 ;
    LAYER V2 ;
      RECT 624 152 656 184 ;
    LAYER V2 ;
      RECT 688 3932 720 3964 ;
    LAYER V2 ;
      RECT 752 152 784 184 ;
    LAYER V2 ;
      RECT 816 3932 848 3964 ;
    LAYER V2 ;
      RECT 880 152 912 184 ;
    LAYER V2 ;
      RECT 944 3932 976 3964 ;
    LAYER V2 ;
      RECT 1008 152 1040 184 ;
    LAYER V2 ;
      RECT 1072 3932 1104 3964 ;
    LAYER V2 ;
      RECT 1136 152 1168 184 ;
    LAYER V2 ;
      RECT 1200 3932 1232 3964 ;
    LAYER V2 ;
      RECT 1264 152 1296 184 ;
    LAYER V2 ;
      RECT 1328 3932 1360 3964 ;
    LAYER V2 ;
      RECT 1392 152 1424 184 ;
    LAYER V2 ;
      RECT 1456 3932 1488 3964 ;
    LAYER V2 ;
      RECT 1520 152 1552 184 ;
    LAYER V2 ;
      RECT 1584 3932 1616 3964 ;
    LAYER V2 ;
      RECT 1648 152 1680 184 ;
    LAYER V2 ;
      RECT 1712 3932 1744 3964 ;
    LAYER V2 ;
      RECT 1776 152 1808 184 ;
    LAYER V2 ;
      RECT 1840 3932 1872 3964 ;
    LAYER V2 ;
      RECT 1904 152 1936 184 ;
    LAYER V2 ;
      RECT 1968 3932 2000 3964 ;
    LAYER V2 ;
      RECT 2032 152 2064 184 ;
    LAYER V2 ;
      RECT 2096 3932 2128 3964 ;
    LAYER V2 ;
      RECT 2160 152 2192 184 ;
    LAYER V2 ;
      RECT 2224 3932 2256 3964 ;
    LAYER V2 ;
      RECT 2288 152 2320 184 ;
    LAYER V2 ;
      RECT 2352 3932 2384 3964 ;
    LAYER V2 ;
      RECT 2416 152 2448 184 ;
    LAYER V2 ;
      RECT 2480 3932 2512 3964 ;
    LAYER V2 ;
      RECT 2544 152 2576 184 ;
    LAYER V2 ;
      RECT 2608 3932 2640 3964 ;
    LAYER V2 ;
      RECT 2672 152 2704 184 ;
    LAYER V2 ;
      RECT 2736 3932 2768 3964 ;
    LAYER V2 ;
      RECT 2800 152 2832 184 ;
    LAYER V2 ;
      RECT 2864 3932 2896 3964 ;
    LAYER V2 ;
      RECT 2928 152 2960 184 ;
    LAYER V2 ;
      RECT 2992 3932 3024 3964 ;
    LAYER V2 ;
      RECT 3056 152 3088 184 ;
    LAYER V2 ;
      RECT 3120 3932 3152 3964 ;
    LAYER V2 ;
      RECT 3184 152 3216 184 ;
    LAYER V2 ;
      RECT 3248 3932 3280 3964 ;
    LAYER V2 ;
      RECT 3312 152 3344 184 ;
    LAYER V2 ;
      RECT 3376 3932 3408 3964 ;
    LAYER V2 ;
      RECT 3440 152 3472 184 ;
    LAYER V2 ;
      RECT 3504 3932 3536 3964 ;
    LAYER V2 ;
      RECT 3568 152 3600 184 ;
    LAYER V2 ;
      RECT 3632 3932 3664 3964 ;
    LAYER V2 ;
      RECT 3696 152 3728 184 ;
    LAYER V2 ;
      RECT 3760 3932 3792 3964 ;
    LAYER V2 ;
      RECT 3824 152 3856 184 ;
    LAYER V2 ;
      RECT 3888 3932 3920 3964 ;
    LAYER V2 ;
      RECT 3952 152 3984 184 ;
    LAYER V2 ;
      RECT 4016 3932 4048 3964 ;
    LAYER V2 ;
      RECT 4144 152 4176 184 ;
    LAYER V2 ;
      RECT 4144 280 4176 312 ;
    LAYER V2 ;
      RECT 4144 408 4176 440 ;
    LAYER V2 ;
      RECT 4144 536 4176 568 ;
    LAYER V2 ;
      RECT 4144 664 4176 696 ;
    LAYER V2 ;
      RECT 4144 792 4176 824 ;
    LAYER V2 ;
      RECT 4144 920 4176 952 ;
    LAYER V2 ;
      RECT 4144 1048 4176 1080 ;
    LAYER V2 ;
      RECT 4144 1176 4176 1208 ;
    LAYER V2 ;
      RECT 4144 1304 4176 1336 ;
    LAYER V2 ;
      RECT 4144 1432 4176 1464 ;
    LAYER V2 ;
      RECT 4144 1560 4176 1592 ;
    LAYER V2 ;
      RECT 4144 1688 4176 1720 ;
    LAYER V2 ;
      RECT 4144 1816 4176 1848 ;
    LAYER V2 ;
      RECT 4144 1944 4176 1976 ;
    LAYER V2 ;
      RECT 4144 2072 4176 2104 ;
    LAYER V2 ;
      RECT 4144 2200 4176 2232 ;
    LAYER V2 ;
      RECT 4144 2328 4176 2360 ;
    LAYER V2 ;
      RECT 4144 2456 4176 2488 ;
    LAYER V2 ;
      RECT 4144 2584 4176 2616 ;
    LAYER V2 ;
      RECT 4144 2712 4176 2744 ;
    LAYER V2 ;
      RECT 4144 2840 4176 2872 ;
    LAYER V2 ;
      RECT 4144 2968 4176 3000 ;
    LAYER V2 ;
      RECT 4144 3096 4176 3128 ;
    LAYER V2 ;
      RECT 4144 3224 4176 3256 ;
    LAYER V2 ;
      RECT 4144 3352 4176 3384 ;
    LAYER V2 ;
      RECT 4144 3480 4176 3512 ;
    LAYER V2 ;
      RECT 4144 3608 4176 3640 ;
    LAYER V2 ;
      RECT 4144 3736 4176 3768 ;
    LAYER V2 ;
      RECT 4144 3864 4176 3896 ;
  END
END CAP_2T_8193393
