MACRO CAP_2T_57809468
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CAP_2T_57809468 0 0 ;
  SIZE 6080 BY 5796 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44 5612 6036 5644 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44 152 6036 184 ;
    END
  END PLUS
  OBS
    LAYER M1 ;
      RECT 304 132 336 5664 ;
    LAYER M1 ;
      RECT 368 132 400 5664 ;
    LAYER M1 ;
      RECT 432 132 464 5664 ;
    LAYER M1 ;
      RECT 496 132 528 5664 ;
    LAYER M1 ;
      RECT 560 132 592 5664 ;
    LAYER M1 ;
      RECT 624 132 656 5664 ;
    LAYER M1 ;
      RECT 688 132 720 5664 ;
    LAYER M1 ;
      RECT 752 132 784 5664 ;
    LAYER M1 ;
      RECT 816 132 848 5664 ;
    LAYER M1 ;
      RECT 880 132 912 5664 ;
    LAYER M1 ;
      RECT 944 132 976 5664 ;
    LAYER M1 ;
      RECT 1008 132 1040 5664 ;
    LAYER M1 ;
      RECT 1072 132 1104 5664 ;
    LAYER M1 ;
      RECT 1136 132 1168 5664 ;
    LAYER M1 ;
      RECT 1200 132 1232 5664 ;
    LAYER M1 ;
      RECT 1264 132 1296 5664 ;
    LAYER M1 ;
      RECT 1328 132 1360 5664 ;
    LAYER M1 ;
      RECT 1392 132 1424 5664 ;
    LAYER M1 ;
      RECT 1456 132 1488 5664 ;
    LAYER M1 ;
      RECT 1520 132 1552 5664 ;
    LAYER M1 ;
      RECT 1584 132 1616 5664 ;
    LAYER M1 ;
      RECT 1648 132 1680 5664 ;
    LAYER M1 ;
      RECT 1712 132 1744 5664 ;
    LAYER M1 ;
      RECT 1776 132 1808 5664 ;
    LAYER M1 ;
      RECT 1840 132 1872 5664 ;
    LAYER M1 ;
      RECT 1904 132 1936 5664 ;
    LAYER M1 ;
      RECT 1968 132 2000 5664 ;
    LAYER M1 ;
      RECT 2032 132 2064 5664 ;
    LAYER M1 ;
      RECT 2096 132 2128 5664 ;
    LAYER M1 ;
      RECT 2160 132 2192 5664 ;
    LAYER M1 ;
      RECT 2224 132 2256 5664 ;
    LAYER M1 ;
      RECT 2288 132 2320 5664 ;
    LAYER M1 ;
      RECT 2352 132 2384 5664 ;
    LAYER M1 ;
      RECT 2416 132 2448 5664 ;
    LAYER M1 ;
      RECT 2480 132 2512 5664 ;
    LAYER M1 ;
      RECT 2544 132 2576 5664 ;
    LAYER M1 ;
      RECT 2608 132 2640 5664 ;
    LAYER M1 ;
      RECT 2672 132 2704 5664 ;
    LAYER M1 ;
      RECT 2736 132 2768 5664 ;
    LAYER M1 ;
      RECT 2800 132 2832 5664 ;
    LAYER M1 ;
      RECT 2864 132 2896 5664 ;
    LAYER M1 ;
      RECT 2928 132 2960 5664 ;
    LAYER M1 ;
      RECT 2992 132 3024 5664 ;
    LAYER M1 ;
      RECT 3056 132 3088 5664 ;
    LAYER M1 ;
      RECT 3120 132 3152 5664 ;
    LAYER M1 ;
      RECT 3184 132 3216 5664 ;
    LAYER M1 ;
      RECT 3248 132 3280 5664 ;
    LAYER M1 ;
      RECT 3312 132 3344 5664 ;
    LAYER M1 ;
      RECT 3376 132 3408 5664 ;
    LAYER M1 ;
      RECT 3440 132 3472 5664 ;
    LAYER M1 ;
      RECT 3504 132 3536 5664 ;
    LAYER M1 ;
      RECT 3568 132 3600 5664 ;
    LAYER M1 ;
      RECT 3632 132 3664 5664 ;
    LAYER M1 ;
      RECT 3696 132 3728 5664 ;
    LAYER M1 ;
      RECT 3760 132 3792 5664 ;
    LAYER M1 ;
      RECT 3824 132 3856 5664 ;
    LAYER M1 ;
      RECT 3888 132 3920 5664 ;
    LAYER M1 ;
      RECT 3952 132 3984 5664 ;
    LAYER M1 ;
      RECT 4016 132 4048 5664 ;
    LAYER M1 ;
      RECT 4080 132 4112 5664 ;
    LAYER M1 ;
      RECT 4144 132 4176 5664 ;
    LAYER M1 ;
      RECT 4208 132 4240 5664 ;
    LAYER M1 ;
      RECT 4272 132 4304 5664 ;
    LAYER M1 ;
      RECT 4336 132 4368 5664 ;
    LAYER M1 ;
      RECT 4400 132 4432 5664 ;
    LAYER M1 ;
      RECT 4464 132 4496 5664 ;
    LAYER M1 ;
      RECT 4528 132 4560 5664 ;
    LAYER M1 ;
      RECT 4592 132 4624 5664 ;
    LAYER M1 ;
      RECT 4656 132 4688 5664 ;
    LAYER M1 ;
      RECT 4720 132 4752 5664 ;
    LAYER M1 ;
      RECT 4784 132 4816 5664 ;
    LAYER M1 ;
      RECT 4848 132 4880 5664 ;
    LAYER M1 ;
      RECT 4912 132 4944 5664 ;
    LAYER M1 ;
      RECT 4976 132 5008 5664 ;
    LAYER M1 ;
      RECT 5040 132 5072 5664 ;
    LAYER M1 ;
      RECT 5104 132 5136 5664 ;
    LAYER M1 ;
      RECT 5168 132 5200 5664 ;
    LAYER M1 ;
      RECT 5232 132 5264 5664 ;
    LAYER M1 ;
      RECT 5296 132 5328 5664 ;
    LAYER M1 ;
      RECT 5360 132 5392 5664 ;
    LAYER M1 ;
      RECT 5424 132 5456 5664 ;
    LAYER M1 ;
      RECT 5488 132 5520 5664 ;
    LAYER M1 ;
      RECT 5552 132 5584 5664 ;
    LAYER M1 ;
      RECT 5616 132 5648 5664 ;
    LAYER M1 ;
      RECT 5680 132 5712 5664 ;
    LAYER M1 ;
      RECT 5744 132 5776 5664 ;
    LAYER M2 ;
      RECT 284 216 5796 248 ;
    LAYER M2 ;
      RECT 284 280 5796 312 ;
    LAYER M2 ;
      RECT 284 344 5796 376 ;
    LAYER M2 ;
      RECT 284 408 5796 440 ;
    LAYER M2 ;
      RECT 284 472 5796 504 ;
    LAYER M2 ;
      RECT 284 536 5796 568 ;
    LAYER M2 ;
      RECT 284 600 5796 632 ;
    LAYER M2 ;
      RECT 284 664 5796 696 ;
    LAYER M2 ;
      RECT 284 728 5796 760 ;
    LAYER M2 ;
      RECT 284 792 5796 824 ;
    LAYER M2 ;
      RECT 284 856 5796 888 ;
    LAYER M2 ;
      RECT 284 920 5796 952 ;
    LAYER M2 ;
      RECT 284 984 5796 1016 ;
    LAYER M2 ;
      RECT 284 1048 5796 1080 ;
    LAYER M2 ;
      RECT 284 1112 5796 1144 ;
    LAYER M2 ;
      RECT 284 1176 5796 1208 ;
    LAYER M2 ;
      RECT 284 1240 5796 1272 ;
    LAYER M2 ;
      RECT 284 1304 5796 1336 ;
    LAYER M2 ;
      RECT 284 1368 5796 1400 ;
    LAYER M2 ;
      RECT 284 1432 5796 1464 ;
    LAYER M2 ;
      RECT 284 1496 5796 1528 ;
    LAYER M2 ;
      RECT 284 1560 5796 1592 ;
    LAYER M2 ;
      RECT 284 1624 5796 1656 ;
    LAYER M2 ;
      RECT 284 1688 5796 1720 ;
    LAYER M2 ;
      RECT 284 1752 5796 1784 ;
    LAYER M2 ;
      RECT 284 1816 5796 1848 ;
    LAYER M2 ;
      RECT 284 1880 5796 1912 ;
    LAYER M2 ;
      RECT 284 1944 5796 1976 ;
    LAYER M2 ;
      RECT 284 2008 5796 2040 ;
    LAYER M2 ;
      RECT 284 2072 5796 2104 ;
    LAYER M2 ;
      RECT 284 2136 5796 2168 ;
    LAYER M2 ;
      RECT 284 2200 5796 2232 ;
    LAYER M2 ;
      RECT 284 2264 5796 2296 ;
    LAYER M2 ;
      RECT 284 2328 5796 2360 ;
    LAYER M2 ;
      RECT 284 2392 5796 2424 ;
    LAYER M2 ;
      RECT 284 2456 5796 2488 ;
    LAYER M2 ;
      RECT 284 2520 5796 2552 ;
    LAYER M2 ;
      RECT 284 2584 5796 2616 ;
    LAYER M2 ;
      RECT 284 2648 5796 2680 ;
    LAYER M2 ;
      RECT 284 2712 5796 2744 ;
    LAYER M2 ;
      RECT 284 2776 5796 2808 ;
    LAYER M2 ;
      RECT 284 2840 5796 2872 ;
    LAYER M2 ;
      RECT 284 2904 5796 2936 ;
    LAYER M2 ;
      RECT 284 2968 5796 3000 ;
    LAYER M2 ;
      RECT 284 3032 5796 3064 ;
    LAYER M2 ;
      RECT 284 3096 5796 3128 ;
    LAYER M2 ;
      RECT 284 3160 5796 3192 ;
    LAYER M2 ;
      RECT 284 3224 5796 3256 ;
    LAYER M2 ;
      RECT 284 3288 5796 3320 ;
    LAYER M2 ;
      RECT 284 3352 5796 3384 ;
    LAYER M2 ;
      RECT 284 3416 5796 3448 ;
    LAYER M2 ;
      RECT 284 3480 5796 3512 ;
    LAYER M2 ;
      RECT 284 3544 5796 3576 ;
    LAYER M2 ;
      RECT 284 3608 5796 3640 ;
    LAYER M2 ;
      RECT 284 3672 5796 3704 ;
    LAYER M2 ;
      RECT 284 3736 5796 3768 ;
    LAYER M2 ;
      RECT 284 3800 5796 3832 ;
    LAYER M2 ;
      RECT 284 3864 5796 3896 ;
    LAYER M2 ;
      RECT 284 3928 5796 3960 ;
    LAYER M2 ;
      RECT 284 3992 5796 4024 ;
    LAYER M2 ;
      RECT 284 4056 5796 4088 ;
    LAYER M2 ;
      RECT 284 4120 5796 4152 ;
    LAYER M2 ;
      RECT 284 4184 5796 4216 ;
    LAYER M2 ;
      RECT 284 4248 5796 4280 ;
    LAYER M2 ;
      RECT 284 4312 5796 4344 ;
    LAYER M2 ;
      RECT 284 4376 5796 4408 ;
    LAYER M2 ;
      RECT 284 4440 5796 4472 ;
    LAYER M2 ;
      RECT 284 4504 5796 4536 ;
    LAYER M2 ;
      RECT 284 4568 5796 4600 ;
    LAYER M2 ;
      RECT 284 4632 5796 4664 ;
    LAYER M2 ;
      RECT 284 4696 5796 4728 ;
    LAYER M2 ;
      RECT 284 4760 5796 4792 ;
    LAYER M2 ;
      RECT 284 4824 5796 4856 ;
    LAYER M2 ;
      RECT 284 4888 5796 4920 ;
    LAYER M2 ;
      RECT 284 4952 5796 4984 ;
    LAYER M2 ;
      RECT 284 5016 5796 5048 ;
    LAYER M2 ;
      RECT 284 5080 5796 5112 ;
    LAYER M2 ;
      RECT 284 5144 5796 5176 ;
    LAYER M2 ;
      RECT 284 5208 5796 5240 ;
    LAYER M2 ;
      RECT 284 5272 5796 5304 ;
    LAYER M2 ;
      RECT 284 5336 5796 5368 ;
    LAYER M2 ;
      RECT 284 5400 5796 5432 ;
    LAYER M2 ;
      RECT 284 5464 5796 5496 ;
    LAYER M2 ;
      RECT 284 5528 5796 5560 ;
    LAYER V1 ;
      RECT 304 216 336 248 ;
    LAYER V1 ;
      RECT 304 344 336 376 ;
    LAYER V1 ;
      RECT 304 472 336 504 ;
    LAYER V1 ;
      RECT 304 600 336 632 ;
    LAYER V1 ;
      RECT 304 728 336 760 ;
    LAYER V1 ;
      RECT 304 856 336 888 ;
    LAYER V1 ;
      RECT 304 984 336 1016 ;
    LAYER V1 ;
      RECT 304 1112 336 1144 ;
    LAYER V1 ;
      RECT 304 1240 336 1272 ;
    LAYER V1 ;
      RECT 304 1368 336 1400 ;
    LAYER V1 ;
      RECT 304 1496 336 1528 ;
    LAYER V1 ;
      RECT 304 1624 336 1656 ;
    LAYER V1 ;
      RECT 304 1752 336 1784 ;
    LAYER V1 ;
      RECT 304 1880 336 1912 ;
    LAYER V1 ;
      RECT 304 2008 336 2040 ;
    LAYER V1 ;
      RECT 304 2136 336 2168 ;
    LAYER V1 ;
      RECT 304 2264 336 2296 ;
    LAYER V1 ;
      RECT 304 2392 336 2424 ;
    LAYER V1 ;
      RECT 304 2520 336 2552 ;
    LAYER V1 ;
      RECT 304 2648 336 2680 ;
    LAYER V1 ;
      RECT 304 2776 336 2808 ;
    LAYER V1 ;
      RECT 304 2904 336 2936 ;
    LAYER V1 ;
      RECT 304 3032 336 3064 ;
    LAYER V1 ;
      RECT 304 3160 336 3192 ;
    LAYER V1 ;
      RECT 304 3288 336 3320 ;
    LAYER V1 ;
      RECT 304 3416 336 3448 ;
    LAYER V1 ;
      RECT 304 3544 336 3576 ;
    LAYER V1 ;
      RECT 304 3672 336 3704 ;
    LAYER V1 ;
      RECT 304 3800 336 3832 ;
    LAYER V1 ;
      RECT 304 3928 336 3960 ;
    LAYER V1 ;
      RECT 304 4056 336 4088 ;
    LAYER V1 ;
      RECT 304 4184 336 4216 ;
    LAYER V1 ;
      RECT 304 4312 336 4344 ;
    LAYER V1 ;
      RECT 304 4440 336 4472 ;
    LAYER V1 ;
      RECT 304 4568 336 4600 ;
    LAYER V1 ;
      RECT 304 4696 336 4728 ;
    LAYER V1 ;
      RECT 304 4824 336 4856 ;
    LAYER V1 ;
      RECT 304 4952 336 4984 ;
    LAYER V1 ;
      RECT 304 5080 336 5112 ;
    LAYER V1 ;
      RECT 304 5208 336 5240 ;
    LAYER V1 ;
      RECT 304 5336 336 5368 ;
    LAYER V1 ;
      RECT 304 5464 336 5496 ;
    LAYER V1 ;
      RECT 304 5612 336 5644 ;
    LAYER V1 ;
      RECT 368 152 400 184 ;
    LAYER V1 ;
      RECT 432 5612 464 5644 ;
    LAYER V1 ;
      RECT 496 152 528 184 ;
    LAYER V1 ;
      RECT 560 5612 592 5644 ;
    LAYER V1 ;
      RECT 624 152 656 184 ;
    LAYER V1 ;
      RECT 688 5612 720 5644 ;
    LAYER V1 ;
      RECT 752 152 784 184 ;
    LAYER V1 ;
      RECT 816 5612 848 5644 ;
    LAYER V1 ;
      RECT 880 152 912 184 ;
    LAYER V1 ;
      RECT 944 5612 976 5644 ;
    LAYER V1 ;
      RECT 1008 152 1040 184 ;
    LAYER V1 ;
      RECT 1072 5612 1104 5644 ;
    LAYER V1 ;
      RECT 1136 152 1168 184 ;
    LAYER V1 ;
      RECT 1200 5612 1232 5644 ;
    LAYER V1 ;
      RECT 1264 152 1296 184 ;
    LAYER V1 ;
      RECT 1328 5612 1360 5644 ;
    LAYER V1 ;
      RECT 1392 152 1424 184 ;
    LAYER V1 ;
      RECT 1456 5612 1488 5644 ;
    LAYER V1 ;
      RECT 1520 152 1552 184 ;
    LAYER V1 ;
      RECT 1584 5612 1616 5644 ;
    LAYER V1 ;
      RECT 1648 152 1680 184 ;
    LAYER V1 ;
      RECT 1712 5612 1744 5644 ;
    LAYER V1 ;
      RECT 1776 152 1808 184 ;
    LAYER V1 ;
      RECT 1840 5612 1872 5644 ;
    LAYER V1 ;
      RECT 1904 152 1936 184 ;
    LAYER V1 ;
      RECT 1968 5612 2000 5644 ;
    LAYER V1 ;
      RECT 2032 152 2064 184 ;
    LAYER V1 ;
      RECT 2096 5612 2128 5644 ;
    LAYER V1 ;
      RECT 2160 152 2192 184 ;
    LAYER V1 ;
      RECT 2224 5612 2256 5644 ;
    LAYER V1 ;
      RECT 2288 152 2320 184 ;
    LAYER V1 ;
      RECT 2352 5612 2384 5644 ;
    LAYER V1 ;
      RECT 2416 152 2448 184 ;
    LAYER V1 ;
      RECT 2480 5612 2512 5644 ;
    LAYER V1 ;
      RECT 2544 152 2576 184 ;
    LAYER V1 ;
      RECT 2608 5612 2640 5644 ;
    LAYER V1 ;
      RECT 2672 152 2704 184 ;
    LAYER V1 ;
      RECT 2736 5612 2768 5644 ;
    LAYER V1 ;
      RECT 2800 152 2832 184 ;
    LAYER V1 ;
      RECT 2864 5612 2896 5644 ;
    LAYER V1 ;
      RECT 2928 152 2960 184 ;
    LAYER V1 ;
      RECT 2992 5612 3024 5644 ;
    LAYER V1 ;
      RECT 3056 152 3088 184 ;
    LAYER V1 ;
      RECT 3120 5612 3152 5644 ;
    LAYER V1 ;
      RECT 3184 152 3216 184 ;
    LAYER V1 ;
      RECT 3248 5612 3280 5644 ;
    LAYER V1 ;
      RECT 3312 152 3344 184 ;
    LAYER V1 ;
      RECT 3376 5612 3408 5644 ;
    LAYER V1 ;
      RECT 3440 152 3472 184 ;
    LAYER V1 ;
      RECT 3504 5612 3536 5644 ;
    LAYER V1 ;
      RECT 3568 152 3600 184 ;
    LAYER V1 ;
      RECT 3632 5612 3664 5644 ;
    LAYER V1 ;
      RECT 3696 152 3728 184 ;
    LAYER V1 ;
      RECT 3760 5612 3792 5644 ;
    LAYER V1 ;
      RECT 3824 152 3856 184 ;
    LAYER V1 ;
      RECT 3888 5612 3920 5644 ;
    LAYER V1 ;
      RECT 3952 152 3984 184 ;
    LAYER V1 ;
      RECT 4016 5612 4048 5644 ;
    LAYER V1 ;
      RECT 4080 152 4112 184 ;
    LAYER V1 ;
      RECT 4144 5612 4176 5644 ;
    LAYER V1 ;
      RECT 4208 152 4240 184 ;
    LAYER V1 ;
      RECT 4272 5612 4304 5644 ;
    LAYER V1 ;
      RECT 4336 152 4368 184 ;
    LAYER V1 ;
      RECT 4400 5612 4432 5644 ;
    LAYER V1 ;
      RECT 4464 152 4496 184 ;
    LAYER V1 ;
      RECT 4528 5612 4560 5644 ;
    LAYER V1 ;
      RECT 4592 152 4624 184 ;
    LAYER V1 ;
      RECT 4656 5612 4688 5644 ;
    LAYER V1 ;
      RECT 4720 152 4752 184 ;
    LAYER V1 ;
      RECT 4784 5612 4816 5644 ;
    LAYER V1 ;
      RECT 4848 152 4880 184 ;
    LAYER V1 ;
      RECT 4912 5612 4944 5644 ;
    LAYER V1 ;
      RECT 4976 152 5008 184 ;
    LAYER V1 ;
      RECT 5040 5612 5072 5644 ;
    LAYER V1 ;
      RECT 5104 152 5136 184 ;
    LAYER V1 ;
      RECT 5168 5612 5200 5644 ;
    LAYER V1 ;
      RECT 5232 152 5264 184 ;
    LAYER V1 ;
      RECT 5296 5612 5328 5644 ;
    LAYER V1 ;
      RECT 5360 152 5392 184 ;
    LAYER V1 ;
      RECT 5424 5612 5456 5644 ;
    LAYER V1 ;
      RECT 5488 152 5520 184 ;
    LAYER V1 ;
      RECT 5552 5612 5584 5644 ;
    LAYER V1 ;
      RECT 5616 152 5648 184 ;
    LAYER V1 ;
      RECT 5680 5612 5712 5644 ;
    LAYER V1 ;
      RECT 5744 152 5776 184 ;
    LAYER V1 ;
      RECT 5744 280 5776 312 ;
    LAYER V1 ;
      RECT 5744 408 5776 440 ;
    LAYER V1 ;
      RECT 5744 536 5776 568 ;
    LAYER V1 ;
      RECT 5744 664 5776 696 ;
    LAYER V1 ;
      RECT 5744 792 5776 824 ;
    LAYER V1 ;
      RECT 5744 920 5776 952 ;
    LAYER V1 ;
      RECT 5744 1048 5776 1080 ;
    LAYER V1 ;
      RECT 5744 1176 5776 1208 ;
    LAYER V1 ;
      RECT 5744 1304 5776 1336 ;
    LAYER V1 ;
      RECT 5744 1432 5776 1464 ;
    LAYER V1 ;
      RECT 5744 1560 5776 1592 ;
    LAYER V1 ;
      RECT 5744 1688 5776 1720 ;
    LAYER V1 ;
      RECT 5744 1816 5776 1848 ;
    LAYER V1 ;
      RECT 5744 1944 5776 1976 ;
    LAYER V1 ;
      RECT 5744 2072 5776 2104 ;
    LAYER V1 ;
      RECT 5744 2200 5776 2232 ;
    LAYER V1 ;
      RECT 5744 2328 5776 2360 ;
    LAYER V1 ;
      RECT 5744 2456 5776 2488 ;
    LAYER V1 ;
      RECT 5744 2584 5776 2616 ;
    LAYER V1 ;
      RECT 5744 2712 5776 2744 ;
    LAYER V1 ;
      RECT 5744 2840 5776 2872 ;
    LAYER V1 ;
      RECT 5744 2968 5776 3000 ;
    LAYER V1 ;
      RECT 5744 3096 5776 3128 ;
    LAYER V1 ;
      RECT 5744 3224 5776 3256 ;
    LAYER V1 ;
      RECT 5744 3352 5776 3384 ;
    LAYER V1 ;
      RECT 5744 3480 5776 3512 ;
    LAYER V1 ;
      RECT 5744 3608 5776 3640 ;
    LAYER V1 ;
      RECT 5744 3736 5776 3768 ;
    LAYER V1 ;
      RECT 5744 3864 5776 3896 ;
    LAYER V1 ;
      RECT 5744 3992 5776 4024 ;
    LAYER V1 ;
      RECT 5744 4120 5776 4152 ;
    LAYER V1 ;
      RECT 5744 4248 5776 4280 ;
    LAYER V1 ;
      RECT 5744 4376 5776 4408 ;
    LAYER V1 ;
      RECT 5744 4504 5776 4536 ;
    LAYER V1 ;
      RECT 5744 4632 5776 4664 ;
    LAYER V1 ;
      RECT 5744 4760 5776 4792 ;
    LAYER V1 ;
      RECT 5744 4888 5776 4920 ;
    LAYER V1 ;
      RECT 5744 5016 5776 5048 ;
    LAYER V1 ;
      RECT 5744 5144 5776 5176 ;
    LAYER V1 ;
      RECT 5744 5272 5776 5304 ;
    LAYER V1 ;
      RECT 5744 5400 5776 5432 ;
    LAYER V1 ;
      RECT 5744 5528 5776 5560 ;
    LAYER M3 ;
      RECT 304 132 336 5664 ;
    LAYER M3 ;
      RECT 368 132 400 5664 ;
    LAYER M3 ;
      RECT 432 132 464 5664 ;
    LAYER M3 ;
      RECT 496 132 528 5664 ;
    LAYER M3 ;
      RECT 560 132 592 5664 ;
    LAYER M3 ;
      RECT 624 132 656 5664 ;
    LAYER M3 ;
      RECT 688 132 720 5664 ;
    LAYER M3 ;
      RECT 752 132 784 5664 ;
    LAYER M3 ;
      RECT 816 132 848 5664 ;
    LAYER M3 ;
      RECT 880 132 912 5664 ;
    LAYER M3 ;
      RECT 944 132 976 5664 ;
    LAYER M3 ;
      RECT 1008 132 1040 5664 ;
    LAYER M3 ;
      RECT 1072 132 1104 5664 ;
    LAYER M3 ;
      RECT 1136 132 1168 5664 ;
    LAYER M3 ;
      RECT 1200 132 1232 5664 ;
    LAYER M3 ;
      RECT 1264 132 1296 5664 ;
    LAYER M3 ;
      RECT 1328 132 1360 5664 ;
    LAYER M3 ;
      RECT 1392 132 1424 5664 ;
    LAYER M3 ;
      RECT 1456 132 1488 5664 ;
    LAYER M3 ;
      RECT 1520 132 1552 5664 ;
    LAYER M3 ;
      RECT 1584 132 1616 5664 ;
    LAYER M3 ;
      RECT 1648 132 1680 5664 ;
    LAYER M3 ;
      RECT 1712 132 1744 5664 ;
    LAYER M3 ;
      RECT 1776 132 1808 5664 ;
    LAYER M3 ;
      RECT 1840 132 1872 5664 ;
    LAYER M3 ;
      RECT 1904 132 1936 5664 ;
    LAYER M3 ;
      RECT 1968 132 2000 5664 ;
    LAYER M3 ;
      RECT 2032 132 2064 5664 ;
    LAYER M3 ;
      RECT 2096 132 2128 5664 ;
    LAYER M3 ;
      RECT 2160 132 2192 5664 ;
    LAYER M3 ;
      RECT 2224 132 2256 5664 ;
    LAYER M3 ;
      RECT 2288 132 2320 5664 ;
    LAYER M3 ;
      RECT 2352 132 2384 5664 ;
    LAYER M3 ;
      RECT 2416 132 2448 5664 ;
    LAYER M3 ;
      RECT 2480 132 2512 5664 ;
    LAYER M3 ;
      RECT 2544 132 2576 5664 ;
    LAYER M3 ;
      RECT 2608 132 2640 5664 ;
    LAYER M3 ;
      RECT 2672 132 2704 5664 ;
    LAYER M3 ;
      RECT 2736 132 2768 5664 ;
    LAYER M3 ;
      RECT 2800 132 2832 5664 ;
    LAYER M3 ;
      RECT 2864 132 2896 5664 ;
    LAYER M3 ;
      RECT 2928 132 2960 5664 ;
    LAYER M3 ;
      RECT 2992 132 3024 5664 ;
    LAYER M3 ;
      RECT 3056 132 3088 5664 ;
    LAYER M3 ;
      RECT 3120 132 3152 5664 ;
    LAYER M3 ;
      RECT 3184 132 3216 5664 ;
    LAYER M3 ;
      RECT 3248 132 3280 5664 ;
    LAYER M3 ;
      RECT 3312 132 3344 5664 ;
    LAYER M3 ;
      RECT 3376 132 3408 5664 ;
    LAYER M3 ;
      RECT 3440 132 3472 5664 ;
    LAYER M3 ;
      RECT 3504 132 3536 5664 ;
    LAYER M3 ;
      RECT 3568 132 3600 5664 ;
    LAYER M3 ;
      RECT 3632 132 3664 5664 ;
    LAYER M3 ;
      RECT 3696 132 3728 5664 ;
    LAYER M3 ;
      RECT 3760 132 3792 5664 ;
    LAYER M3 ;
      RECT 3824 132 3856 5664 ;
    LAYER M3 ;
      RECT 3888 132 3920 5664 ;
    LAYER M3 ;
      RECT 3952 132 3984 5664 ;
    LAYER M3 ;
      RECT 4016 132 4048 5664 ;
    LAYER M3 ;
      RECT 4080 132 4112 5664 ;
    LAYER M3 ;
      RECT 4144 132 4176 5664 ;
    LAYER M3 ;
      RECT 4208 132 4240 5664 ;
    LAYER M3 ;
      RECT 4272 132 4304 5664 ;
    LAYER M3 ;
      RECT 4336 132 4368 5664 ;
    LAYER M3 ;
      RECT 4400 132 4432 5664 ;
    LAYER M3 ;
      RECT 4464 132 4496 5664 ;
    LAYER M3 ;
      RECT 4528 132 4560 5664 ;
    LAYER M3 ;
      RECT 4592 132 4624 5664 ;
    LAYER M3 ;
      RECT 4656 132 4688 5664 ;
    LAYER M3 ;
      RECT 4720 132 4752 5664 ;
    LAYER M3 ;
      RECT 4784 132 4816 5664 ;
    LAYER M3 ;
      RECT 4848 132 4880 5664 ;
    LAYER M3 ;
      RECT 4912 132 4944 5664 ;
    LAYER M3 ;
      RECT 4976 132 5008 5664 ;
    LAYER M3 ;
      RECT 5040 132 5072 5664 ;
    LAYER M3 ;
      RECT 5104 132 5136 5664 ;
    LAYER M3 ;
      RECT 5168 132 5200 5664 ;
    LAYER M3 ;
      RECT 5232 132 5264 5664 ;
    LAYER M3 ;
      RECT 5296 132 5328 5664 ;
    LAYER M3 ;
      RECT 5360 132 5392 5664 ;
    LAYER M3 ;
      RECT 5424 132 5456 5664 ;
    LAYER M3 ;
      RECT 5488 132 5520 5664 ;
    LAYER M3 ;
      RECT 5552 132 5584 5664 ;
    LAYER M3 ;
      RECT 5616 132 5648 5664 ;
    LAYER M3 ;
      RECT 5680 132 5712 5664 ;
    LAYER M3 ;
      RECT 5740 132 5780 5664 ;
    LAYER V2 ;
      RECT 304 216 336 248 ;
    LAYER V2 ;
      RECT 304 344 336 376 ;
    LAYER V2 ;
      RECT 304 472 336 504 ;
    LAYER V2 ;
      RECT 304 600 336 632 ;
    LAYER V2 ;
      RECT 304 728 336 760 ;
    LAYER V2 ;
      RECT 304 856 336 888 ;
    LAYER V2 ;
      RECT 304 984 336 1016 ;
    LAYER V2 ;
      RECT 304 1112 336 1144 ;
    LAYER V2 ;
      RECT 304 1240 336 1272 ;
    LAYER V2 ;
      RECT 304 1368 336 1400 ;
    LAYER V2 ;
      RECT 304 1496 336 1528 ;
    LAYER V2 ;
      RECT 304 1624 336 1656 ;
    LAYER V2 ;
      RECT 304 1752 336 1784 ;
    LAYER V2 ;
      RECT 304 1880 336 1912 ;
    LAYER V2 ;
      RECT 304 2008 336 2040 ;
    LAYER V2 ;
      RECT 304 2136 336 2168 ;
    LAYER V2 ;
      RECT 304 2264 336 2296 ;
    LAYER V2 ;
      RECT 304 2392 336 2424 ;
    LAYER V2 ;
      RECT 304 2520 336 2552 ;
    LAYER V2 ;
      RECT 304 2648 336 2680 ;
    LAYER V2 ;
      RECT 304 2776 336 2808 ;
    LAYER V2 ;
      RECT 304 2904 336 2936 ;
    LAYER V2 ;
      RECT 304 3032 336 3064 ;
    LAYER V2 ;
      RECT 304 3160 336 3192 ;
    LAYER V2 ;
      RECT 304 3288 336 3320 ;
    LAYER V2 ;
      RECT 304 3416 336 3448 ;
    LAYER V2 ;
      RECT 304 3544 336 3576 ;
    LAYER V2 ;
      RECT 304 3672 336 3704 ;
    LAYER V2 ;
      RECT 304 3800 336 3832 ;
    LAYER V2 ;
      RECT 304 3928 336 3960 ;
    LAYER V2 ;
      RECT 304 4056 336 4088 ;
    LAYER V2 ;
      RECT 304 4184 336 4216 ;
    LAYER V2 ;
      RECT 304 4312 336 4344 ;
    LAYER V2 ;
      RECT 304 4440 336 4472 ;
    LAYER V2 ;
      RECT 304 4568 336 4600 ;
    LAYER V2 ;
      RECT 304 4696 336 4728 ;
    LAYER V2 ;
      RECT 304 4824 336 4856 ;
    LAYER V2 ;
      RECT 304 4952 336 4984 ;
    LAYER V2 ;
      RECT 304 5080 336 5112 ;
    LAYER V2 ;
      RECT 304 5208 336 5240 ;
    LAYER V2 ;
      RECT 304 5336 336 5368 ;
    LAYER V2 ;
      RECT 304 5464 336 5496 ;
    LAYER V2 ;
      RECT 304 5612 336 5644 ;
    LAYER V2 ;
      RECT 368 152 400 184 ;
    LAYER V2 ;
      RECT 432 5612 464 5644 ;
    LAYER V2 ;
      RECT 496 152 528 184 ;
    LAYER V2 ;
      RECT 560 5612 592 5644 ;
    LAYER V2 ;
      RECT 624 152 656 184 ;
    LAYER V2 ;
      RECT 688 5612 720 5644 ;
    LAYER V2 ;
      RECT 752 152 784 184 ;
    LAYER V2 ;
      RECT 816 5612 848 5644 ;
    LAYER V2 ;
      RECT 880 152 912 184 ;
    LAYER V2 ;
      RECT 944 5612 976 5644 ;
    LAYER V2 ;
      RECT 1008 152 1040 184 ;
    LAYER V2 ;
      RECT 1072 5612 1104 5644 ;
    LAYER V2 ;
      RECT 1136 152 1168 184 ;
    LAYER V2 ;
      RECT 1200 5612 1232 5644 ;
    LAYER V2 ;
      RECT 1264 152 1296 184 ;
    LAYER V2 ;
      RECT 1328 5612 1360 5644 ;
    LAYER V2 ;
      RECT 1392 152 1424 184 ;
    LAYER V2 ;
      RECT 1456 5612 1488 5644 ;
    LAYER V2 ;
      RECT 1520 152 1552 184 ;
    LAYER V2 ;
      RECT 1584 5612 1616 5644 ;
    LAYER V2 ;
      RECT 1648 152 1680 184 ;
    LAYER V2 ;
      RECT 1712 5612 1744 5644 ;
    LAYER V2 ;
      RECT 1776 152 1808 184 ;
    LAYER V2 ;
      RECT 1840 5612 1872 5644 ;
    LAYER V2 ;
      RECT 1904 152 1936 184 ;
    LAYER V2 ;
      RECT 1968 5612 2000 5644 ;
    LAYER V2 ;
      RECT 2032 152 2064 184 ;
    LAYER V2 ;
      RECT 2096 5612 2128 5644 ;
    LAYER V2 ;
      RECT 2160 152 2192 184 ;
    LAYER V2 ;
      RECT 2224 5612 2256 5644 ;
    LAYER V2 ;
      RECT 2288 152 2320 184 ;
    LAYER V2 ;
      RECT 2352 5612 2384 5644 ;
    LAYER V2 ;
      RECT 2416 152 2448 184 ;
    LAYER V2 ;
      RECT 2480 5612 2512 5644 ;
    LAYER V2 ;
      RECT 2544 152 2576 184 ;
    LAYER V2 ;
      RECT 2608 5612 2640 5644 ;
    LAYER V2 ;
      RECT 2672 152 2704 184 ;
    LAYER V2 ;
      RECT 2736 5612 2768 5644 ;
    LAYER V2 ;
      RECT 2800 152 2832 184 ;
    LAYER V2 ;
      RECT 2864 5612 2896 5644 ;
    LAYER V2 ;
      RECT 2928 152 2960 184 ;
    LAYER V2 ;
      RECT 2992 5612 3024 5644 ;
    LAYER V2 ;
      RECT 3056 152 3088 184 ;
    LAYER V2 ;
      RECT 3120 5612 3152 5644 ;
    LAYER V2 ;
      RECT 3184 152 3216 184 ;
    LAYER V2 ;
      RECT 3248 5612 3280 5644 ;
    LAYER V2 ;
      RECT 3312 152 3344 184 ;
    LAYER V2 ;
      RECT 3376 5612 3408 5644 ;
    LAYER V2 ;
      RECT 3440 152 3472 184 ;
    LAYER V2 ;
      RECT 3504 5612 3536 5644 ;
    LAYER V2 ;
      RECT 3568 152 3600 184 ;
    LAYER V2 ;
      RECT 3632 5612 3664 5644 ;
    LAYER V2 ;
      RECT 3696 152 3728 184 ;
    LAYER V2 ;
      RECT 3760 5612 3792 5644 ;
    LAYER V2 ;
      RECT 3824 152 3856 184 ;
    LAYER V2 ;
      RECT 3888 5612 3920 5644 ;
    LAYER V2 ;
      RECT 3952 152 3984 184 ;
    LAYER V2 ;
      RECT 4016 5612 4048 5644 ;
    LAYER V2 ;
      RECT 4080 152 4112 184 ;
    LAYER V2 ;
      RECT 4144 5612 4176 5644 ;
    LAYER V2 ;
      RECT 4208 152 4240 184 ;
    LAYER V2 ;
      RECT 4272 5612 4304 5644 ;
    LAYER V2 ;
      RECT 4336 152 4368 184 ;
    LAYER V2 ;
      RECT 4400 5612 4432 5644 ;
    LAYER V2 ;
      RECT 4464 152 4496 184 ;
    LAYER V2 ;
      RECT 4528 5612 4560 5644 ;
    LAYER V2 ;
      RECT 4592 152 4624 184 ;
    LAYER V2 ;
      RECT 4656 5612 4688 5644 ;
    LAYER V2 ;
      RECT 4720 152 4752 184 ;
    LAYER V2 ;
      RECT 4784 5612 4816 5644 ;
    LAYER V2 ;
      RECT 4848 152 4880 184 ;
    LAYER V2 ;
      RECT 4912 5612 4944 5644 ;
    LAYER V2 ;
      RECT 4976 152 5008 184 ;
    LAYER V2 ;
      RECT 5040 5612 5072 5644 ;
    LAYER V2 ;
      RECT 5104 152 5136 184 ;
    LAYER V2 ;
      RECT 5168 5612 5200 5644 ;
    LAYER V2 ;
      RECT 5232 152 5264 184 ;
    LAYER V2 ;
      RECT 5296 5612 5328 5644 ;
    LAYER V2 ;
      RECT 5360 152 5392 184 ;
    LAYER V2 ;
      RECT 5424 5612 5456 5644 ;
    LAYER V2 ;
      RECT 5488 152 5520 184 ;
    LAYER V2 ;
      RECT 5552 5612 5584 5644 ;
    LAYER V2 ;
      RECT 5616 152 5648 184 ;
    LAYER V2 ;
      RECT 5680 5612 5712 5644 ;
    LAYER V2 ;
      RECT 5744 152 5776 184 ;
    LAYER V2 ;
      RECT 5744 280 5776 312 ;
    LAYER V2 ;
      RECT 5744 408 5776 440 ;
    LAYER V2 ;
      RECT 5744 536 5776 568 ;
    LAYER V2 ;
      RECT 5744 664 5776 696 ;
    LAYER V2 ;
      RECT 5744 792 5776 824 ;
    LAYER V2 ;
      RECT 5744 920 5776 952 ;
    LAYER V2 ;
      RECT 5744 1048 5776 1080 ;
    LAYER V2 ;
      RECT 5744 1176 5776 1208 ;
    LAYER V2 ;
      RECT 5744 1304 5776 1336 ;
    LAYER V2 ;
      RECT 5744 1432 5776 1464 ;
    LAYER V2 ;
      RECT 5744 1560 5776 1592 ;
    LAYER V2 ;
      RECT 5744 1688 5776 1720 ;
    LAYER V2 ;
      RECT 5744 1816 5776 1848 ;
    LAYER V2 ;
      RECT 5744 1944 5776 1976 ;
    LAYER V2 ;
      RECT 5744 2072 5776 2104 ;
    LAYER V2 ;
      RECT 5744 2200 5776 2232 ;
    LAYER V2 ;
      RECT 5744 2328 5776 2360 ;
    LAYER V2 ;
      RECT 5744 2456 5776 2488 ;
    LAYER V2 ;
      RECT 5744 2584 5776 2616 ;
    LAYER V2 ;
      RECT 5744 2712 5776 2744 ;
    LAYER V2 ;
      RECT 5744 2840 5776 2872 ;
    LAYER V2 ;
      RECT 5744 2968 5776 3000 ;
    LAYER V2 ;
      RECT 5744 3096 5776 3128 ;
    LAYER V2 ;
      RECT 5744 3224 5776 3256 ;
    LAYER V2 ;
      RECT 5744 3352 5776 3384 ;
    LAYER V2 ;
      RECT 5744 3480 5776 3512 ;
    LAYER V2 ;
      RECT 5744 3608 5776 3640 ;
    LAYER V2 ;
      RECT 5744 3736 5776 3768 ;
    LAYER V2 ;
      RECT 5744 3864 5776 3896 ;
    LAYER V2 ;
      RECT 5744 3992 5776 4024 ;
    LAYER V2 ;
      RECT 5744 4120 5776 4152 ;
    LAYER V2 ;
      RECT 5744 4248 5776 4280 ;
    LAYER V2 ;
      RECT 5744 4376 5776 4408 ;
    LAYER V2 ;
      RECT 5744 4504 5776 4536 ;
    LAYER V2 ;
      RECT 5744 4632 5776 4664 ;
    LAYER V2 ;
      RECT 5744 4760 5776 4792 ;
    LAYER V2 ;
      RECT 5744 4888 5776 4920 ;
    LAYER V2 ;
      RECT 5744 5016 5776 5048 ;
    LAYER V2 ;
      RECT 5744 5144 5776 5176 ;
    LAYER V2 ;
      RECT 5744 5272 5776 5304 ;
    LAYER V2 ;
      RECT 5744 5400 5776 5432 ;
    LAYER V2 ;
      RECT 5744 5528 5776 5560 ;
  END
END CAP_2T_57809468
