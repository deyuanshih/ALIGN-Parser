MACRO CMC_S_NMOS_B_2722902_X2_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CMC_S_NMOS_B_2722902_X2_Y1 0 0 ;
  SIZE 2560 BY 2352 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 1748 2276 1780 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 68 996 100 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1564 152 2276 184 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 908 2276 940 ;
    END
  END G
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204 236 1076 268 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1484 320 2356 352 ;
    END
  END SB
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1644 336 1884 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 944 48 976 792 ;
    LAYER M1 ;
      RECT 944 888 976 1128 ;
    LAYER M1 ;
      RECT 944 1644 976 1884 ;
    LAYER M1 ;
      RECT 864 48 896 792 ;
    LAYER M1 ;
      RECT 1024 48 1056 792 ;
    LAYER M1 ;
      RECT 1584 48 1616 792 ;
    LAYER M1 ;
      RECT 1584 888 1616 1128 ;
    LAYER M1 ;
      RECT 1584 1644 1616 1884 ;
    LAYER M1 ;
      RECT 1504 48 1536 792 ;
    LAYER M1 ;
      RECT 1664 48 1696 792 ;
    LAYER M1 ;
      RECT 2224 48 2256 792 ;
    LAYER M1 ;
      RECT 2224 888 2256 1128 ;
    LAYER M1 ;
      RECT 2224 1644 2256 1884 ;
    LAYER M1 ;
      RECT 2144 48 2176 792 ;
    LAYER M1 ;
      RECT 2304 48 2336 792 ;
    LAYER V1 ;
      RECT 944 68 976 100 ;
    LAYER V1 ;
      RECT 944 908 976 940 ;
    LAYER V1 ;
      RECT 944 1748 976 1780 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1748 336 1780 ;
    LAYER V1 ;
      RECT 2224 152 2256 184 ;
    LAYER V1 ;
      RECT 2224 908 2256 940 ;
    LAYER V1 ;
      RECT 2224 1748 2256 1780 ;
    LAYER V1 ;
      RECT 1584 152 1616 184 ;
    LAYER V1 ;
      RECT 1584 908 1616 940 ;
    LAYER V1 ;
      RECT 1584 1748 1616 1780 ;
    LAYER V1 ;
      RECT 864 236 896 268 ;
    LAYER V1 ;
      RECT 1024 236 1056 268 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 2144 320 2176 352 ;
    LAYER V1 ;
      RECT 1664 320 1696 352 ;
    LAYER V1 ;
      RECT 1504 320 1536 352 ;
    LAYER V1 ;
      RECT 2304 320 2336 352 ;
    LAYER V0 ;
      RECT 304 398 336 430 ;
    LAYER V0 ;
      RECT 304 482 336 514 ;
    LAYER V0 ;
      RECT 304 566 336 598 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1748 336 1780 ;
    LAYER V0 ;
      RECT 224 398 256 430 ;
    LAYER V0 ;
      RECT 224 482 256 514 ;
    LAYER V0 ;
      RECT 224 566 256 598 ;
    LAYER V0 ;
      RECT 384 398 416 430 ;
    LAYER V0 ;
      RECT 384 482 416 514 ;
    LAYER V0 ;
      RECT 384 566 416 598 ;
    LAYER V0 ;
      RECT 944 398 976 430 ;
    LAYER V0 ;
      RECT 944 482 976 514 ;
    LAYER V0 ;
      RECT 944 566 976 598 ;
    LAYER V0 ;
      RECT 944 908 976 940 ;
    LAYER V0 ;
      RECT 944 1748 976 1780 ;
    LAYER V0 ;
      RECT 864 398 896 430 ;
    LAYER V0 ;
      RECT 864 482 896 514 ;
    LAYER V0 ;
      RECT 864 566 896 598 ;
    LAYER V0 ;
      RECT 1024 398 1056 430 ;
    LAYER V0 ;
      RECT 1024 482 1056 514 ;
    LAYER V0 ;
      RECT 1024 566 1056 598 ;
    LAYER V0 ;
      RECT 1584 398 1616 430 ;
    LAYER V0 ;
      RECT 1584 482 1616 514 ;
    LAYER V0 ;
      RECT 1584 566 1616 598 ;
    LAYER V0 ;
      RECT 1584 908 1616 940 ;
    LAYER V0 ;
      RECT 1584 1748 1616 1780 ;
    LAYER V0 ;
      RECT 1504 398 1536 430 ;
    LAYER V0 ;
      RECT 1504 482 1536 514 ;
    LAYER V0 ;
      RECT 1504 566 1536 598 ;
    LAYER V0 ;
      RECT 1664 398 1696 430 ;
    LAYER V0 ;
      RECT 1664 482 1696 514 ;
    LAYER V0 ;
      RECT 1664 566 1696 598 ;
    LAYER V0 ;
      RECT 2224 398 2256 430 ;
    LAYER V0 ;
      RECT 2224 482 2256 514 ;
    LAYER V0 ;
      RECT 2224 566 2256 598 ;
    LAYER V0 ;
      RECT 2224 908 2256 940 ;
    LAYER V0 ;
      RECT 2224 1748 2256 1780 ;
    LAYER V0 ;
      RECT 2144 398 2176 430 ;
    LAYER V0 ;
      RECT 2144 482 2176 514 ;
    LAYER V0 ;
      RECT 2144 566 2176 598 ;
    LAYER V0 ;
      RECT 2304 398 2336 430 ;
    LAYER V0 ;
      RECT 2304 482 2336 514 ;
    LAYER V0 ;
      RECT 2304 566 2336 598 ;
  END
END CMC_S_NMOS_B_2722902_X2_Y1
