MACRO DP_NMOS_B_40344802_X1_Y3
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_40344802_X1_Y3 0 0 ;
  SIZE 800 BY 4704 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 4100 516 4132 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 60 48 100 2472 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 140 132 180 2556 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 220 888 260 3312 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 300 972 340 3396 ;
    END
  END GB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 380 216 420 2640 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1224 336 1968 ;
    LAYER M1 ;
      RECT 304 2064 336 2304 ;
    LAYER M1 ;
      RECT 304 2400 336 3144 ;
    LAYER M1 ;
      RECT 304 3240 336 3480 ;
    LAYER M1 ;
      RECT 304 3996 336 4236 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 224 1224 256 1968 ;
    LAYER M1 ;
      RECT 224 2400 256 3144 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 384 1224 416 1968 ;
    LAYER M1 ;
      RECT 384 2400 416 3144 ;
    LAYER M1 ;
      RECT 464 48 496 792 ;
    LAYER M1 ;
      RECT 464 888 496 1128 ;
    LAYER M1 ;
      RECT 464 1224 496 1968 ;
    LAYER M1 ;
      RECT 464 2064 496 2304 ;
    LAYER M1 ;
      RECT 464 2400 496 3144 ;
    LAYER M1 ;
      RECT 464 3240 496 3480 ;
    LAYER M1 ;
      RECT 464 3996 496 4236 ;
    LAYER M1 ;
      RECT 544 48 576 792 ;
    LAYER M1 ;
      RECT 544 1224 576 1968 ;
    LAYER M1 ;
      RECT 544 2400 576 3144 ;
    LAYER M2 ;
      RECT 44 68 356 100 ;
    LAYER M2 ;
      RECT 124 152 516 184 ;
    LAYER M2 ;
      RECT 124 908 356 940 ;
    LAYER M2 ;
      RECT 284 992 516 1024 ;
    LAYER M2 ;
      RECT 204 236 596 268 ;
    LAYER M2 ;
      RECT 44 1244 516 1276 ;
    LAYER M2 ;
      RECT 124 1328 356 1360 ;
    LAYER M2 ;
      RECT 204 2084 516 2116 ;
    LAYER M2 ;
      RECT 124 2168 356 2200 ;
    LAYER M2 ;
      RECT 204 1412 596 1444 ;
    LAYER M2 ;
      RECT 44 2420 356 2452 ;
    LAYER M2 ;
      RECT 124 2504 516 2536 ;
    LAYER M2 ;
      RECT 124 3260 356 3292 ;
    LAYER M2 ;
      RECT 284 3344 516 3376 ;
    LAYER M2 ;
      RECT 204 2588 596 2620 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1328 336 1360 ;
    LAYER V1 ;
      RECT 304 2168 336 2200 ;
    LAYER V1 ;
      RECT 304 2420 336 2452 ;
    LAYER V1 ;
      RECT 304 3260 336 3292 ;
    LAYER V1 ;
      RECT 304 4100 336 4132 ;
    LAYER V1 ;
      RECT 464 152 496 184 ;
    LAYER V1 ;
      RECT 464 992 496 1024 ;
    LAYER V1 ;
      RECT 464 1244 496 1276 ;
    LAYER V1 ;
      RECT 464 2084 496 2116 ;
    LAYER V1 ;
      RECT 464 2504 496 2536 ;
    LAYER V1 ;
      RECT 464 3344 496 3376 ;
    LAYER V1 ;
      RECT 464 4100 496 4132 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 224 1412 256 1444 ;
    LAYER V1 ;
      RECT 224 2588 256 2620 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 384 1412 416 1444 ;
    LAYER V1 ;
      RECT 384 2588 416 2620 ;
    LAYER V1 ;
      RECT 544 236 576 268 ;
    LAYER V1 ;
      RECT 544 1412 576 1444 ;
    LAYER V1 ;
      RECT 544 2588 576 2620 ;
    LAYER V2 ;
      RECT 64 68 96 100 ;
    LAYER V2 ;
      RECT 64 1244 96 1276 ;
    LAYER V2 ;
      RECT 64 2420 96 2452 ;
    LAYER V2 ;
      RECT 144 152 176 184 ;
    LAYER V2 ;
      RECT 144 1328 176 1360 ;
    LAYER V2 ;
      RECT 144 2504 176 2536 ;
    LAYER V2 ;
      RECT 224 908 256 940 ;
    LAYER V2 ;
      RECT 224 2084 256 2116 ;
    LAYER V2 ;
      RECT 224 3260 256 3292 ;
    LAYER V2 ;
      RECT 304 992 336 1024 ;
    LAYER V2 ;
      RECT 304 2168 336 2200 ;
    LAYER V2 ;
      RECT 304 3344 336 3376 ;
    LAYER V2 ;
      RECT 384 236 416 268 ;
    LAYER V2 ;
      RECT 384 1412 416 1444 ;
    LAYER V2 ;
      RECT 384 2588 416 2620 ;
    LAYER V0 ;
      RECT 304 335 336 367 ;
    LAYER V0 ;
      RECT 304 419 336 451 ;
    LAYER V0 ;
      RECT 304 503 336 535 ;
    LAYER V0 ;
      RECT 304 587 336 619 ;
    LAYER V0 ;
      RECT 304 671 336 703 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1511 336 1543 ;
    LAYER V0 ;
      RECT 304 1595 336 1627 ;
    LAYER V0 ;
      RECT 304 1679 336 1711 ;
    LAYER V0 ;
      RECT 304 1763 336 1795 ;
    LAYER V0 ;
      RECT 304 1847 336 1879 ;
    LAYER V0 ;
      RECT 304 2084 336 2116 ;
    LAYER V0 ;
      RECT 304 2687 336 2719 ;
    LAYER V0 ;
      RECT 304 2771 336 2803 ;
    LAYER V0 ;
      RECT 304 2855 336 2887 ;
    LAYER V0 ;
      RECT 304 2939 336 2971 ;
    LAYER V0 ;
      RECT 304 3023 336 3055 ;
    LAYER V0 ;
      RECT 304 3260 336 3292 ;
    LAYER V0 ;
      RECT 304 4100 336 4132 ;
    LAYER V0 ;
      RECT 304 4100 336 4132 ;
    LAYER V0 ;
      RECT 304 4100 336 4132 ;
    LAYER V0 ;
      RECT 224 335 256 367 ;
    LAYER V0 ;
      RECT 224 419 256 451 ;
    LAYER V0 ;
      RECT 224 503 256 535 ;
    LAYER V0 ;
      RECT 224 587 256 619 ;
    LAYER V0 ;
      RECT 224 671 256 703 ;
    LAYER V0 ;
      RECT 224 1511 256 1543 ;
    LAYER V0 ;
      RECT 224 1595 256 1627 ;
    LAYER V0 ;
      RECT 224 1679 256 1711 ;
    LAYER V0 ;
      RECT 224 1763 256 1795 ;
    LAYER V0 ;
      RECT 224 1847 256 1879 ;
    LAYER V0 ;
      RECT 224 2687 256 2719 ;
    LAYER V0 ;
      RECT 224 2771 256 2803 ;
    LAYER V0 ;
      RECT 224 2855 256 2887 ;
    LAYER V0 ;
      RECT 224 2939 256 2971 ;
    LAYER V0 ;
      RECT 224 3023 256 3055 ;
    LAYER V0 ;
      RECT 384 335 416 367 ;
    LAYER V0 ;
      RECT 384 335 416 367 ;
    LAYER V0 ;
      RECT 384 419 416 451 ;
    LAYER V0 ;
      RECT 384 419 416 451 ;
    LAYER V0 ;
      RECT 384 503 416 535 ;
    LAYER V0 ;
      RECT 384 503 416 535 ;
    LAYER V0 ;
      RECT 384 587 416 619 ;
    LAYER V0 ;
      RECT 384 587 416 619 ;
    LAYER V0 ;
      RECT 384 671 416 703 ;
    LAYER V0 ;
      RECT 384 671 416 703 ;
    LAYER V0 ;
      RECT 384 1511 416 1543 ;
    LAYER V0 ;
      RECT 384 1511 416 1543 ;
    LAYER V0 ;
      RECT 384 1595 416 1627 ;
    LAYER V0 ;
      RECT 384 1595 416 1627 ;
    LAYER V0 ;
      RECT 384 1679 416 1711 ;
    LAYER V0 ;
      RECT 384 1679 416 1711 ;
    LAYER V0 ;
      RECT 384 1763 416 1795 ;
    LAYER V0 ;
      RECT 384 1763 416 1795 ;
    LAYER V0 ;
      RECT 384 1847 416 1879 ;
    LAYER V0 ;
      RECT 384 1847 416 1879 ;
    LAYER V0 ;
      RECT 384 2687 416 2719 ;
    LAYER V0 ;
      RECT 384 2687 416 2719 ;
    LAYER V0 ;
      RECT 384 2771 416 2803 ;
    LAYER V0 ;
      RECT 384 2771 416 2803 ;
    LAYER V0 ;
      RECT 384 2855 416 2887 ;
    LAYER V0 ;
      RECT 384 2855 416 2887 ;
    LAYER V0 ;
      RECT 384 2939 416 2971 ;
    LAYER V0 ;
      RECT 384 2939 416 2971 ;
    LAYER V0 ;
      RECT 384 3023 416 3055 ;
    LAYER V0 ;
      RECT 384 3023 416 3055 ;
    LAYER V0 ;
      RECT 464 335 496 367 ;
    LAYER V0 ;
      RECT 464 419 496 451 ;
    LAYER V0 ;
      RECT 464 503 496 535 ;
    LAYER V0 ;
      RECT 464 587 496 619 ;
    LAYER V0 ;
      RECT 464 671 496 703 ;
    LAYER V0 ;
      RECT 464 908 496 940 ;
    LAYER V0 ;
      RECT 464 1511 496 1543 ;
    LAYER V0 ;
      RECT 464 1595 496 1627 ;
    LAYER V0 ;
      RECT 464 1679 496 1711 ;
    LAYER V0 ;
      RECT 464 1763 496 1795 ;
    LAYER V0 ;
      RECT 464 1847 496 1879 ;
    LAYER V0 ;
      RECT 464 2084 496 2116 ;
    LAYER V0 ;
      RECT 464 2687 496 2719 ;
    LAYER V0 ;
      RECT 464 2771 496 2803 ;
    LAYER V0 ;
      RECT 464 2855 496 2887 ;
    LAYER V0 ;
      RECT 464 2939 496 2971 ;
    LAYER V0 ;
      RECT 464 3023 496 3055 ;
    LAYER V0 ;
      RECT 464 3260 496 3292 ;
    LAYER V0 ;
      RECT 464 4100 496 4132 ;
    LAYER V0 ;
      RECT 464 4100 496 4132 ;
    LAYER V0 ;
      RECT 464 4100 496 4132 ;
    LAYER V0 ;
      RECT 544 335 576 367 ;
    LAYER V0 ;
      RECT 544 419 576 451 ;
    LAYER V0 ;
      RECT 544 503 576 535 ;
    LAYER V0 ;
      RECT 544 587 576 619 ;
    LAYER V0 ;
      RECT 544 671 576 703 ;
    LAYER V0 ;
      RECT 544 1511 576 1543 ;
    LAYER V0 ;
      RECT 544 1595 576 1627 ;
    LAYER V0 ;
      RECT 544 1679 576 1711 ;
    LAYER V0 ;
      RECT 544 1763 576 1795 ;
    LAYER V0 ;
      RECT 544 1847 576 1879 ;
    LAYER V0 ;
      RECT 544 2687 576 2719 ;
    LAYER V0 ;
      RECT 544 2771 576 2803 ;
    LAYER V0 ;
      RECT 544 2855 576 2887 ;
    LAYER V0 ;
      RECT 544 2939 576 2971 ;
    LAYER V0 ;
      RECT 544 3023 576 3055 ;
  END
END DP_NMOS_B_40344802_X1_Y3
