.subckt DFCND4BWP_LVT D CP CDN Q QN VDD VSS
MI14_3  net175 net149 VDD VDD plvt w=102.5n l=40n nf=8 nfin=8
MI22_3  Q net149 VDD VDD plvt w=102.5n l=40n nf=8 nfin=8
MI28_3  QN net175 VDD VDD plvt w=102.5n l=40n nf=8 nfin=8
MI23_3  QN net175 VDD VDD plvt w=102.5n l=40n nf=8 nfin=8
MI43  net12 net145 VDD VDD plvt w=30.0n l=40n nf=8 nfin=8
MI39_3  net95 net11 VDD VDD plvt w=102.5n l=40n nf=8 nfin=8
MI6  net9 D net1 VDD plvt w=85n l=40n nf=8 nfin=8
MI26_3  QN net175 VDD VDD plvt w=102.5n l=40n nf=8 nfin=8
MI29_3  QN net175 VDD VDD plvt w=102.5n l=40n nf=8 nfin=8
MI31_3  net11 CP VDD VDD plvt w=102.5n l=40n nf=8 nfin=8
MI27_3  Q net149 VDD VDD plvt w=102.5n l=40n nf=8 nfin=8
MI36_2  net149 CDN VDD VDD plvt w=102.5n l=40n nf=8 nfin=8
MI44  net12 CDN VDD VDD plvt w=30.0n l=40n nf=8 nfin=8
MI17  net175 net95 net24 VDD plvt w=30.0n l=40n nf=8 nfin=8
MI36_1  net149 net24 VDD VDD plvt w=102.5n l=40n nf=8 nfin=8
MI13_3  net145 net9 VDD VDD plvt w=45n l=40n nf=8 nfin=8
MI24_3  Q net149 VDD VDD plvt w=102.5n l=40n nf=8 nfin=8
MI16  net145 net11 net24 VDD plvt w=45n l=40n nf=8 nfin=8
MI30_1  net149 net24 VDD VDD plvt w=70n l=40n nf=8 nfin=8
MI30_2  net149 CDN VDD VDD plvt w=70n l=40n nf=8 nfin=8
MI45  net9 net11 net12 VDD plvt w=30.0n l=40n nf=8 nfin=8
MI25_3  Q net149 VDD VDD plvt w=102.5n l=40n nf=8 nfin=8
MI7  net1 net95 VDD VDD plvt w=85.0n l=40n nf=8 nfin=8
MI26_2  QN net175 VSS VSS nlvt w=77.5n l=40n nf=8 nfin=8
MI24_2  Q net149 VSS VSS nlvt w=77.5n l=40n nf=8 nfin=8
MI29_2  QN net175 VSS VSS nlvt w=77.5n l=40n nf=8 nfin=8
MI30_4  net169 CDN VSS VSS nlvt w=50n l=40n nf=8 nfin=8
MI4  net128 net11 VSS VSS nlvt w=77.5n l=40n nf=8 nfin=8
MI23_2  QN net175 VSS VSS nlvt w=77.5n l=40n nf=8 nfin=8
MI18  net175 net11 net24 VSS nlvt w=30.0n l=40n nf=8 nfin=8
MI13_2  net145 net9 VSS VSS nlvt w=37.5n l=40n nf=8 nfin=8
MI30_3  net149 net24 net169 VSS nlvt w=50n l=40n nf=8 nfin=8
MI15  net145 net95 net24 VSS nlvt w=37.5n l=40n nf=8 nfin=8
MI14_2  net175 net149 VSS VSS nlvt w=47.5n l=40n nf=8 nfin=8
MI25_2  Q net149 VSS VSS nlvt w=77.5n l=40n nf=8 nfin=8
MI39_2  net95 net11 VSS VSS nlvt w=77.5n l=40n nf=8 nfin=8
MI36_3  net149 net24 net132 VSS nlvt w=50n l=40n nf=8 nfin=8
MI5  net9 D net128 VSS nlvt w=77.5n l=40n nf=8 nfin=8
MI31_2  net11 CP VSS VSS nlvt w=77.5n l=40n nf=8 nfin=8
MI49  net112 CDN VSS VSS nlvt w=30.0n l=40n nf=8 nfin=8
MI36_4  net132 CDN VSS VSS nlvt w=50n l=40n nf=8 nfin=8
MI48  net96 net145 net112 VSS nlvt w=30.0n l=40n nf=8 nfin=8
MI27_2  Q net149 VSS VSS nlvt w=77.5n l=40n nf=8 nfin=8
MI28_2  QN net175 VSS VSS nlvt w=77.5n l=40n nf=8 nfin=8
MI22_2  Q net149 VSS VSS nlvt w=77.5n l=40n nf=8 nfin=8
MI47  net9 net95 net96 VSS nlvt w=30.0n l=40n nf=8 nfin=8
.ends DFCND4BWP_LVT