MACRO PMOS_S_32343612_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN PMOS_S_32343612_X1_Y1 0 0 ;
  SIZE 640 BY 2352 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124 68 356 100 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124 908 356 940 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 220 132 260 1800 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1644 336 1884 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M2 ;
      RECT 124 1748 356 1780 ;
    LAYER M2 ;
      RECT 204 152 436 184 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1748 336 1780 ;
    LAYER V1 ;
      RECT 224 152 256 184 ;
    LAYER V1 ;
      RECT 384 152 416 184 ;
    LAYER V2 ;
      RECT 224 152 256 184 ;
    LAYER V2 ;
      RECT 224 1748 256 1780 ;
    LAYER V0 ;
      RECT 304 545 336 577 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1748 336 1780 ;
    LAYER V0 ;
      RECT 224 545 256 577 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
  END
END PMOS_S_32343612_X1_Y1
