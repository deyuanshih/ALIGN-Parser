MACRO CCP_NMOS_23282412_X1_Y4
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CCP_NMOS_23282412_X1_Y4 0 0 ;
  SIZE 800 BY 5880 ;
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 140 48 180 4488 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 220 132 260 4572 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 300 216 340 5328 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1224 336 1968 ;
    LAYER M1 ;
      RECT 304 2064 336 2304 ;
    LAYER M1 ;
      RECT 304 2400 336 3144 ;
    LAYER M1 ;
      RECT 304 3240 336 3480 ;
    LAYER M1 ;
      RECT 304 3576 336 4320 ;
    LAYER M1 ;
      RECT 304 4416 336 4656 ;
    LAYER M1 ;
      RECT 304 5172 336 5412 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 224 1224 256 1968 ;
    LAYER M1 ;
      RECT 224 2400 256 3144 ;
    LAYER M1 ;
      RECT 224 3576 256 4320 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 384 1224 416 1968 ;
    LAYER M1 ;
      RECT 384 2400 416 3144 ;
    LAYER M1 ;
      RECT 384 3576 416 4320 ;
    LAYER M1 ;
      RECT 464 48 496 792 ;
    LAYER M1 ;
      RECT 464 888 496 1128 ;
    LAYER M1 ;
      RECT 464 1224 496 1968 ;
    LAYER M1 ;
      RECT 464 2064 496 2304 ;
    LAYER M1 ;
      RECT 464 2400 496 3144 ;
    LAYER M1 ;
      RECT 464 3240 496 3480 ;
    LAYER M1 ;
      RECT 464 3576 496 4320 ;
    LAYER M1 ;
      RECT 464 4416 496 4656 ;
    LAYER M1 ;
      RECT 464 5172 496 5412 ;
    LAYER M1 ;
      RECT 544 48 576 792 ;
    LAYER M1 ;
      RECT 544 1224 576 1968 ;
    LAYER M1 ;
      RECT 544 2400 576 3144 ;
    LAYER M1 ;
      RECT 544 3576 576 4320 ;
    LAYER M2 ;
      RECT 124 908 516 940 ;
    LAYER M2 ;
      RECT 124 68 356 100 ;
    LAYER M2 ;
      RECT 124 992 356 1024 ;
    LAYER M2 ;
      RECT 204 152 516 184 ;
    LAYER M2 ;
      RECT 204 236 596 268 ;
    LAYER M2 ;
      RECT 124 2084 356 2116 ;
    LAYER M2 ;
      RECT 124 1244 516 1276 ;
    LAYER M2 ;
      RECT 204 2168 516 2200 ;
    LAYER M2 ;
      RECT 124 1328 356 1360 ;
    LAYER M2 ;
      RECT 204 1412 596 1444 ;
    LAYER M2 ;
      RECT 124 3260 516 3292 ;
    LAYER M2 ;
      RECT 124 2420 356 2452 ;
    LAYER M2 ;
      RECT 124 3344 356 3376 ;
    LAYER M2 ;
      RECT 204 2504 516 2536 ;
    LAYER M2 ;
      RECT 204 2588 596 2620 ;
    LAYER M2 ;
      RECT 124 4436 356 4468 ;
    LAYER M2 ;
      RECT 124 3596 516 3628 ;
    LAYER M2 ;
      RECT 204 4520 516 4552 ;
    LAYER M2 ;
      RECT 124 3680 356 3712 ;
    LAYER M2 ;
      RECT 284 5276 516 5308 ;
    LAYER M2 ;
      RECT 204 3764 596 3796 ;
    LAYER V1 ;
      RECT 464 152 496 184 ;
    LAYER V1 ;
      RECT 464 908 496 940 ;
    LAYER V1 ;
      RECT 464 1244 496 1276 ;
    LAYER V1 ;
      RECT 464 2168 496 2200 ;
    LAYER V1 ;
      RECT 464 2504 496 2536 ;
    LAYER V1 ;
      RECT 464 3260 496 3292 ;
    LAYER V1 ;
      RECT 464 3596 496 3628 ;
    LAYER V1 ;
      RECT 464 4520 496 4552 ;
    LAYER V1 ;
      RECT 464 5276 496 5308 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 992 336 1024 ;
    LAYER V1 ;
      RECT 304 1328 336 1360 ;
    LAYER V1 ;
      RECT 304 2084 336 2116 ;
    LAYER V1 ;
      RECT 304 2420 336 2452 ;
    LAYER V1 ;
      RECT 304 3344 336 3376 ;
    LAYER V1 ;
      RECT 304 3680 336 3712 ;
    LAYER V1 ;
      RECT 304 4436 336 4468 ;
    LAYER V1 ;
      RECT 304 5276 336 5308 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 224 1412 256 1444 ;
    LAYER V1 ;
      RECT 224 2588 256 2620 ;
    LAYER V1 ;
      RECT 224 3764 256 3796 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 384 1412 416 1444 ;
    LAYER V1 ;
      RECT 384 2588 416 2620 ;
    LAYER V1 ;
      RECT 384 3764 416 3796 ;
    LAYER V1 ;
      RECT 544 236 576 268 ;
    LAYER V1 ;
      RECT 544 1412 576 1444 ;
    LAYER V1 ;
      RECT 544 2588 576 2620 ;
    LAYER V1 ;
      RECT 544 3764 576 3796 ;
    LAYER V2 ;
      RECT 144 68 176 100 ;
    LAYER V2 ;
      RECT 144 908 176 940 ;
    LAYER V2 ;
      RECT 144 1244 176 1276 ;
    LAYER V2 ;
      RECT 144 2084 176 2116 ;
    LAYER V2 ;
      RECT 144 2420 176 2452 ;
    LAYER V2 ;
      RECT 144 3260 176 3292 ;
    LAYER V2 ;
      RECT 144 3596 176 3628 ;
    LAYER V2 ;
      RECT 144 4436 176 4468 ;
    LAYER V2 ;
      RECT 224 152 256 184 ;
    LAYER V2 ;
      RECT 224 992 256 1024 ;
    LAYER V2 ;
      RECT 224 1328 256 1360 ;
    LAYER V2 ;
      RECT 224 2168 256 2200 ;
    LAYER V2 ;
      RECT 224 2504 256 2536 ;
    LAYER V2 ;
      RECT 224 3344 256 3376 ;
    LAYER V2 ;
      RECT 224 3680 256 3712 ;
    LAYER V2 ;
      RECT 224 4520 256 4552 ;
    LAYER V2 ;
      RECT 304 236 336 268 ;
    LAYER V2 ;
      RECT 304 1412 336 1444 ;
    LAYER V2 ;
      RECT 304 2588 336 2620 ;
    LAYER V2 ;
      RECT 304 3764 336 3796 ;
    LAYER V2 ;
      RECT 304 5276 336 5308 ;
    LAYER V0 ;
      RECT 304 545 336 577 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1721 336 1753 ;
    LAYER V0 ;
      RECT 304 2084 336 2116 ;
    LAYER V0 ;
      RECT 304 2897 336 2929 ;
    LAYER V0 ;
      RECT 304 3260 336 3292 ;
    LAYER V0 ;
      RECT 304 4073 336 4105 ;
    LAYER V0 ;
      RECT 304 4436 336 4468 ;
    LAYER V0 ;
      RECT 304 5276 336 5308 ;
    LAYER V0 ;
      RECT 304 5276 336 5308 ;
    LAYER V0 ;
      RECT 304 5276 336 5308 ;
    LAYER V0 ;
      RECT 304 5276 336 5308 ;
    LAYER V0 ;
      RECT 224 545 256 577 ;
    LAYER V0 ;
      RECT 224 1721 256 1753 ;
    LAYER V0 ;
      RECT 224 2897 256 2929 ;
    LAYER V0 ;
      RECT 224 4073 256 4105 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 384 1721 416 1753 ;
    LAYER V0 ;
      RECT 384 1721 416 1753 ;
    LAYER V0 ;
      RECT 384 2897 416 2929 ;
    LAYER V0 ;
      RECT 384 2897 416 2929 ;
    LAYER V0 ;
      RECT 384 4073 416 4105 ;
    LAYER V0 ;
      RECT 384 4073 416 4105 ;
    LAYER V0 ;
      RECT 464 545 496 577 ;
    LAYER V0 ;
      RECT 464 908 496 940 ;
    LAYER V0 ;
      RECT 464 1721 496 1753 ;
    LAYER V0 ;
      RECT 464 2084 496 2116 ;
    LAYER V0 ;
      RECT 464 2897 496 2929 ;
    LAYER V0 ;
      RECT 464 3260 496 3292 ;
    LAYER V0 ;
      RECT 464 4073 496 4105 ;
    LAYER V0 ;
      RECT 464 4436 496 4468 ;
    LAYER V0 ;
      RECT 464 5276 496 5308 ;
    LAYER V0 ;
      RECT 464 5276 496 5308 ;
    LAYER V0 ;
      RECT 464 5276 496 5308 ;
    LAYER V0 ;
      RECT 464 5276 496 5308 ;
    LAYER V0 ;
      RECT 544 545 576 577 ;
    LAYER V0 ;
      RECT 544 1721 576 1753 ;
    LAYER V0 ;
      RECT 544 2897 576 2929 ;
    LAYER V0 ;
      RECT 544 4073 576 4105 ;
  END
END CCP_NMOS_23282412_X1_Y4
