MACRO CMC_PMOS_95878848_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_95878848_X1_Y1 0 0 ;
  SIZE 800 BY 2352 ;
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124 68 356 100 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 152 516 184 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 908 516 940 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 380 216 420 1800 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1644 336 1884 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 464 48 496 792 ;
    LAYER M1 ;
      RECT 464 888 496 1128 ;
    LAYER M1 ;
      RECT 464 1644 496 1884 ;
    LAYER M1 ;
      RECT 544 48 576 792 ;
    LAYER M2 ;
      RECT 284 1748 516 1780 ;
    LAYER M2 ;
      RECT 204 236 596 268 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1748 336 1780 ;
    LAYER V1 ;
      RECT 464 152 496 184 ;
    LAYER V1 ;
      RECT 464 908 496 940 ;
    LAYER V1 ;
      RECT 464 1748 496 1780 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 544 236 576 268 ;
    LAYER V2 ;
      RECT 384 236 416 268 ;
    LAYER V2 ;
      RECT 384 1748 416 1780 ;
    LAYER V0 ;
      RECT 304 461 336 493 ;
    LAYER V0 ;
      RECT 304 545 336 577 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1748 336 1780 ;
    LAYER V0 ;
      RECT 224 461 256 493 ;
    LAYER V0 ;
      RECT 224 545 256 577 ;
    LAYER V0 ;
      RECT 384 461 416 493 ;
    LAYER V0 ;
      RECT 384 461 416 493 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 464 461 496 493 ;
    LAYER V0 ;
      RECT 464 545 496 577 ;
    LAYER V0 ;
      RECT 464 908 496 940 ;
    LAYER V0 ;
      RECT 464 1748 496 1780 ;
    LAYER V0 ;
      RECT 544 461 576 493 ;
    LAYER V0 ;
      RECT 544 545 576 577 ;
  END
END CMC_PMOS_95878848_X1_Y1
