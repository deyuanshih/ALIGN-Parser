MACRO SWITCHED_CAPACITOR_FILTER
  ORIGIN 0 0 ;
  FOREIGN SWITCHED_CAPACITOR_FILTER 0 0 ;
  SIZE 58.612 BY 40.204 ;
  PIN ID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 29.5 23.484 29.54 24.396 ;
    END
  END ID
  PIN VBIASN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 29.42 14.244 29.46 15.492 ;
    END
  END VBIASN
  PIN VBIASP1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 29.164 19.64 29.396 19.672 ;
    END
  END VBIASP1
  PIN VBIASP2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 29.404 17.288 29.636 17.32 ;
      LAYER M2 ;
        RECT 28.924 17.288 29.156 17.32 ;
      LAYER M2 ;
        RECT 29.12 17.288 29.44 17.32 ;
    END
  END VBIASP2
  PIN VOUTN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 29.404 16.448 29.636 16.48 ;
      LAYER M3 ;
        RECT 29.18 15 29.22 16.248 ;
      LAYER M2 ;
        RECT 29.36 16.448 29.44 16.48 ;
      LAYER M3 ;
        RECT 29.34 16.359 29.38 16.569 ;
      LAYER M4 ;
        RECT 29.2 16.444 29.36 16.484 ;
      LAYER M3 ;
        RECT 29.18 16.212 29.22 16.464 ;
      LAYER M1 ;
        RECT 58.304 13.068 58.336 13.14 ;
      LAYER M2 ;
        RECT 58.284 13.088 58.356 13.12 ;
      LAYER M1 ;
        RECT 30.704 13.068 30.736 13.14 ;
      LAYER M2 ;
        RECT 30.684 13.088 30.756 13.12 ;
      LAYER M2 ;
        RECT 30.72 13.088 58.32 13.12 ;
      LAYER M2 ;
        RECT 29.404 12.752 29.636 12.784 ;
      LAYER M2 ;
        RECT 30.364 10.316 36.356 10.348 ;
      LAYER M3 ;
        RECT 29.18 13.104 29.22 15.036 ;
      LAYER M2 ;
        RECT 29.2 13.088 30.72 13.12 ;
      LAYER M2 ;
        RECT 29.484 13.088 29.556 13.12 ;
      LAYER M3 ;
        RECT 29.5 12.768 29.54 13.104 ;
      LAYER M2 ;
        RECT 29.484 12.752 29.556 12.784 ;
      LAYER M2 ;
        RECT 36.124 13.088 36.196 13.12 ;
      LAYER M1 ;
        RECT 36.144 10.332 36.176 13.104 ;
      LAYER M2 ;
        RECT 36.124 10.316 36.196 10.348 ;
    END
  END VOUTN
  PIN VOUTP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 28.924 16.448 29.156 16.48 ;
      LAYER M3 ;
        RECT 29.1 15.084 29.14 16.332 ;
      LAYER M2 ;
        RECT 29.084 16.448 29.156 16.48 ;
      LAYER M3 ;
        RECT 29.1 16.296 29.14 16.464 ;
      LAYER M1 ;
        RECT 0.224 13.068 0.256 13.14 ;
      LAYER M2 ;
        RECT 0.204 13.088 0.276 13.12 ;
      LAYER M1 ;
        RECT 27.824 13.068 27.856 13.14 ;
      LAYER M2 ;
        RECT 27.804 13.088 27.876 13.12 ;
      LAYER M2 ;
        RECT 0.24 13.088 27.84 13.12 ;
      LAYER M2 ;
        RECT 28.924 12.668 29.156 12.7 ;
      LAYER M2 ;
        RECT 22.204 10.316 28.196 10.348 ;
      LAYER M3 ;
        RECT 29.1 14.196 29.14 15.12 ;
      LAYER M2 ;
        RECT 28.98 14.18 29.18 14.212 ;
      LAYER M1 ;
        RECT 29.024 13.104 29.056 14.196 ;
      LAYER M2 ;
        RECT 27.84 13.088 29.04 13.12 ;
      LAYER M2 ;
        RECT 29.004 13.088 29.076 13.12 ;
      LAYER M3 ;
        RECT 29.02 12.684 29.06 13.104 ;
      LAYER M2 ;
        RECT 29.004 12.668 29.076 12.7 ;
      LAYER M2 ;
        RECT 27.964 13.088 28.036 13.12 ;
      LAYER M1 ;
        RECT 27.984 10.332 28.016 13.104 ;
      LAYER M2 ;
        RECT 27.964 10.316 28.036 10.348 ;
    END
  END VOUTP
  PIN PHI2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 29.164 5.696 29.396 5.728 ;
      LAYER M2 ;
        RECT 28.204 13.76 28.436 13.792 ;
      LAYER M2 ;
        RECT 30.124 13.76 30.356 13.792 ;
      LAYER M2 ;
        RECT 29.804 6.116 30.036 6.148 ;
      LAYER M2 ;
        RECT 28.524 6.116 28.756 6.148 ;
      LAYER M2 ;
        RECT 29.12 5.696 29.2 5.728 ;
      LAYER M3 ;
        RECT 29.1 5.712 29.14 13.776 ;
      LAYER M2 ;
        RECT 28.4 13.76 29.12 13.792 ;
      LAYER M3 ;
        RECT 29.1 13.736 29.14 13.816 ;
      LAYER M4 ;
        RECT 29.12 13.756 29.28 13.796 ;
      LAYER M3 ;
        RECT 29.26 13.671 29.3 13.881 ;
      LAYER M2 ;
        RECT 29.28 13.76 30.16 13.792 ;
      LAYER M3 ;
        RECT 29.1 6.092 29.14 6.172 ;
      LAYER M2 ;
        RECT 29.12 6.116 29.84 6.148 ;
      LAYER M3 ;
        RECT 29.1 6.092 29.14 6.172 ;
      LAYER M4 ;
        RECT 28.88 6.112 29.12 6.152 ;
      LAYER M3 ;
        RECT 28.86 6.027 28.9 6.237 ;
      LAYER M2 ;
        RECT 28.72 6.116 28.88 6.148 ;
    END
  END PHI2
  PIN AGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 29.084 5.024 29.476 5.056 ;
      LAYER M2 ;
        RECT 28.204 12.92 28.436 12.952 ;
      LAYER M2 ;
        RECT 30.124 12.92 30.356 12.952 ;
      LAYER M2 ;
        RECT 29.804 6.956 30.036 6.988 ;
      LAYER M2 ;
        RECT 28.524 6.956 28.756 6.988 ;
      LAYER M2 ;
        RECT 28.8 5.024 29.12 5.056 ;
      LAYER M1 ;
        RECT 28.784 5.04 28.816 12.936 ;
      LAYER M2 ;
        RECT 28.4 12.92 28.8 12.952 ;
      LAYER M2 ;
        RECT 28.8 12.92 30.16 12.952 ;
      LAYER M1 ;
        RECT 28.784 6.852 28.816 6.924 ;
      LAYER M2 ;
        RECT 28.8 6.872 29 6.904 ;
      LAYER M1 ;
        RECT 28.864 6.84 28.896 7.02 ;
      LAYER M2 ;
        RECT 28.88 6.956 29.84 6.988 ;
      LAYER M2 ;
        RECT 28.72 6.956 28.88 6.988 ;
    END
  END AGND
  PIN PHI1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 28.924 11.912 29.636 11.944 ;
      LAYER M2 ;
        RECT 28.924 1.412 29.636 1.444 ;
      LAYER M2 ;
        RECT 28.924 3.764 29.636 3.796 ;
      LAYER M2 ;
        RECT 29.244 11.912 29.316 11.944 ;
      LAYER M3 ;
        RECT 29.26 1.428 29.3 11.928 ;
      LAYER M2 ;
        RECT 29.244 1.412 29.316 1.444 ;
      LAYER M3 ;
        RECT 29.26 3.74 29.3 3.82 ;
      LAYER M2 ;
        RECT 29.244 3.764 29.316 3.796 ;
    END
  END PHI1
  PIN VINP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 29.484 4.436 29.716 4.468 ;
      LAYER M2 ;
        RECT 36.444 4.856 42.436 4.888 ;
      LAYER M2 ;
        RECT 29.68 4.436 36.48 4.468 ;
      LAYER M1 ;
        RECT 36.464 4.452 36.496 4.872 ;
      LAYER M2 ;
        RECT 36.444 4.856 36.516 4.888 ;
    END
  END VINP
  PIN VINN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 28.844 4.352 29.076 4.384 ;
      LAYER M2 ;
        RECT 16.124 4.856 22.116 4.888 ;
      LAYER M2 ;
        RECT 22.08 4.352 28.88 4.384 ;
      LAYER M1 ;
        RECT 22.064 4.368 22.096 4.872 ;
      LAYER M2 ;
        RECT 22.044 4.856 22.116 4.888 ;
    END
  END VINN
  OBS 
  LAYER M2 ;
        RECT 29.004 22.076 29.716 22.108 ;
  LAYER M1 ;
        RECT 0.064 39.864 0.096 39.936 ;
  LAYER M2 ;
        RECT 0.044 39.884 0.116 39.916 ;
  LAYER M1 ;
        RECT 27.664 39.864 27.696 39.936 ;
  LAYER M2 ;
        RECT 27.644 39.884 27.716 39.916 ;
  LAYER M2 ;
        RECT 0.08 39.884 27.68 39.916 ;
  LAYER M2 ;
        RECT 28.924 2.252 29.156 2.284 ;
  LAYER M2 ;
        RECT 16.124 10.316 22.116 10.348 ;
  LAYER M2 ;
        RECT 29.004 22.076 29.076 22.108 ;
  LAYER M3 ;
        RECT 29.02 22.092 29.06 39.9 ;
  LAYER M2 ;
        RECT 27.68 39.884 29.04 39.916 ;
  LAYER M3 ;
        RECT 29.02 22.052 29.06 22.132 ;
  LAYER M4 ;
        RECT 28.93 22.072 29.07 22.112 ;
  LAYER M3 ;
        RECT 28.94 2.268 28.98 22.092 ;
  LAYER M2 ;
        RECT 28.924 2.252 28.996 2.284 ;
  LAYER M3 ;
        RECT 28.94 10.292 28.98 10.372 ;
  LAYER M4 ;
        RECT 22.08 10.312 28.96 10.352 ;
  LAYER M3 ;
        RECT 22.06 10.227 22.1 10.437 ;
  LAYER M2 ;
        RECT 22.044 10.316 22.116 10.348 ;
  LAYER M2 ;
        RECT 29.004 22.076 29.076 22.108 ;
  LAYER M3 ;
        RECT 29.02 22.056 29.06 22.128 ;
  LAYER M2 ;
        RECT 29.004 39.884 29.076 39.916 ;
  LAYER M3 ;
        RECT 29.02 39.864 29.06 39.936 ;
  LAYER M2 ;
        RECT 29.004 22.076 29.076 22.108 ;
  LAYER M3 ;
        RECT 29.02 22.056 29.06 22.128 ;
  LAYER M2 ;
        RECT 29.004 39.884 29.076 39.916 ;
  LAYER M3 ;
        RECT 29.02 39.864 29.06 39.936 ;
  LAYER M2 ;
        RECT 28.924 2.252 28.996 2.284 ;
  LAYER M3 ;
        RECT 28.94 2.232 28.98 2.304 ;
  LAYER M2 ;
        RECT 29.004 22.076 29.076 22.108 ;
  LAYER M3 ;
        RECT 29.02 22.056 29.06 22.128 ;
  LAYER M2 ;
        RECT 29.004 39.884 29.076 39.916 ;
  LAYER M3 ;
        RECT 29.02 39.864 29.06 39.936 ;
  LAYER M3 ;
        RECT 28.94 22.052 28.98 22.132 ;
  LAYER M4 ;
        RECT 28.92 22.072 29 22.112 ;
  LAYER M3 ;
        RECT 29.02 22.052 29.06 22.132 ;
  LAYER M4 ;
        RECT 29 22.072 29.08 22.112 ;
  LAYER M2 ;
        RECT 28.924 2.252 28.996 2.284 ;
  LAYER M3 ;
        RECT 28.94 2.232 28.98 2.304 ;
  LAYER M2 ;
        RECT 29.004 22.076 29.076 22.108 ;
  LAYER M3 ;
        RECT 29.02 22.056 29.06 22.128 ;
  LAYER M2 ;
        RECT 29.004 39.884 29.076 39.916 ;
  LAYER M3 ;
        RECT 29.02 39.864 29.06 39.936 ;
  LAYER M2 ;
        RECT 22.044 10.316 22.116 10.348 ;
  LAYER M3 ;
        RECT 22.06 10.296 22.1 10.368 ;
  LAYER M2 ;
        RECT 28.924 2.252 28.996 2.284 ;
  LAYER M3 ;
        RECT 28.94 2.232 28.98 2.304 ;
  LAYER M2 ;
        RECT 29.004 22.076 29.076 22.108 ;
  LAYER M3 ;
        RECT 29.02 22.056 29.06 22.128 ;
  LAYER M2 ;
        RECT 29.004 39.884 29.076 39.916 ;
  LAYER M3 ;
        RECT 29.02 39.864 29.06 39.936 ;
  LAYER M3 ;
        RECT 22.06 10.292 22.1 10.372 ;
  LAYER M4 ;
        RECT 22.04 10.312 22.12 10.352 ;
  LAYER M3 ;
        RECT 28.94 10.292 28.98 10.372 ;
  LAYER M4 ;
        RECT 28.92 10.312 29 10.352 ;
  LAYER M2 ;
        RECT 28.924 2.252 28.996 2.284 ;
  LAYER M3 ;
        RECT 28.94 2.232 28.98 2.304 ;
  LAYER M2 ;
        RECT 29.004 22.076 29.076 22.108 ;
  LAYER M3 ;
        RECT 29.02 22.056 29.06 22.128 ;
  LAYER M2 ;
        RECT 29.004 39.884 29.076 39.916 ;
  LAYER M3 ;
        RECT 29.02 39.864 29.06 39.936 ;
  LAYER M3 ;
        RECT 28.94 10.292 28.98 10.372 ;
  LAYER M4 ;
        RECT 28.92 10.312 29 10.352 ;
  LAYER M2 ;
        RECT 28.844 21.992 29.556 22.024 ;
  LAYER M1 ;
        RECT 58.464 39.864 58.496 39.936 ;
  LAYER M2 ;
        RECT 58.444 39.884 58.516 39.916 ;
  LAYER M1 ;
        RECT 30.864 39.864 30.896 39.936 ;
  LAYER M2 ;
        RECT 30.844 39.884 30.916 39.916 ;
  LAYER M2 ;
        RECT 30.88 39.884 58.48 39.916 ;
  LAYER M2 ;
        RECT 29.404 2.168 29.636 2.2 ;
  LAYER M2 ;
        RECT 36.444 10.316 42.436 10.348 ;
  LAYER M2 ;
        RECT 29.52 21.992 29.6 22.024 ;
  LAYER M3 ;
        RECT 29.58 22.008 29.62 39.9 ;
  LAYER M2 ;
        RECT 29.6 39.884 30.88 39.916 ;
  LAYER M3 ;
        RECT 29.58 2.184 29.62 22.008 ;
  LAYER M2 ;
        RECT 29.564 2.168 29.636 2.2 ;
  LAYER M3 ;
        RECT 29.58 10.292 29.62 10.372 ;
  LAYER M4 ;
        RECT 29.6 10.312 36.48 10.352 ;
  LAYER M3 ;
        RECT 36.46 10.227 36.5 10.437 ;
  LAYER M2 ;
        RECT 36.444 10.316 36.516 10.348 ;
  LAYER M2 ;
        RECT 29.564 21.992 29.636 22.024 ;
  LAYER M3 ;
        RECT 29.58 21.972 29.62 22.044 ;
  LAYER M2 ;
        RECT 29.564 39.884 29.636 39.916 ;
  LAYER M3 ;
        RECT 29.58 39.864 29.62 39.936 ;
  LAYER M2 ;
        RECT 29.564 21.992 29.636 22.024 ;
  LAYER M3 ;
        RECT 29.58 21.972 29.62 22.044 ;
  LAYER M2 ;
        RECT 29.564 39.884 29.636 39.916 ;
  LAYER M3 ;
        RECT 29.58 39.864 29.62 39.936 ;
  LAYER M2 ;
        RECT 29.564 2.168 29.636 2.2 ;
  LAYER M3 ;
        RECT 29.58 2.148 29.62 2.22 ;
  LAYER M2 ;
        RECT 29.564 21.992 29.636 22.024 ;
  LAYER M3 ;
        RECT 29.58 21.972 29.62 22.044 ;
  LAYER M2 ;
        RECT 29.564 39.884 29.636 39.916 ;
  LAYER M3 ;
        RECT 29.58 39.864 29.62 39.936 ;
  LAYER M2 ;
        RECT 29.564 2.168 29.636 2.2 ;
  LAYER M3 ;
        RECT 29.58 2.148 29.62 2.22 ;
  LAYER M2 ;
        RECT 29.564 21.992 29.636 22.024 ;
  LAYER M3 ;
        RECT 29.58 21.972 29.62 22.044 ;
  LAYER M2 ;
        RECT 29.564 39.884 29.636 39.916 ;
  LAYER M3 ;
        RECT 29.58 39.864 29.62 39.936 ;
  LAYER M2 ;
        RECT 29.564 2.168 29.636 2.2 ;
  LAYER M3 ;
        RECT 29.58 2.148 29.62 2.22 ;
  LAYER M2 ;
        RECT 29.564 21.992 29.636 22.024 ;
  LAYER M3 ;
        RECT 29.58 21.972 29.62 22.044 ;
  LAYER M2 ;
        RECT 29.564 39.884 29.636 39.916 ;
  LAYER M3 ;
        RECT 29.58 39.864 29.62 39.936 ;
  LAYER M2 ;
        RECT 36.444 10.316 36.516 10.348 ;
  LAYER M3 ;
        RECT 36.46 10.296 36.5 10.368 ;
  LAYER M3 ;
        RECT 29.58 10.292 29.62 10.372 ;
  LAYER M4 ;
        RECT 29.56 10.312 29.64 10.352 ;
  LAYER M3 ;
        RECT 36.46 10.292 36.5 10.372 ;
  LAYER M4 ;
        RECT 36.44 10.312 36.52 10.352 ;
  LAYER M2 ;
        RECT 29.564 2.168 29.636 2.2 ;
  LAYER M3 ;
        RECT 29.58 2.148 29.62 2.22 ;
  LAYER M2 ;
        RECT 29.564 21.992 29.636 22.024 ;
  LAYER M3 ;
        RECT 29.58 21.972 29.62 22.044 ;
  LAYER M2 ;
        RECT 29.564 39.884 29.636 39.916 ;
  LAYER M3 ;
        RECT 29.58 39.864 29.62 39.936 ;
  LAYER M3 ;
        RECT 29.58 10.292 29.62 10.372 ;
  LAYER M4 ;
        RECT 29.56 10.312 29.64 10.352 ;
  LAYER M1 ;
        RECT 48.944 13.236 48.976 13.308 ;
  LAYER M2 ;
        RECT 48.924 13.256 48.996 13.288 ;
  LAYER M1 ;
        RECT 39.744 13.236 39.776 13.308 ;
  LAYER M2 ;
        RECT 39.724 13.256 39.796 13.288 ;
  LAYER M2 ;
        RECT 39.76 13.256 48.96 13.288 ;
  LAYER M2 ;
        RECT 29.484 12.584 29.716 12.616 ;
  LAYER M2 ;
        RECT 30.204 13.004 30.436 13.036 ;
  LAYER M1 ;
        RECT 39.744 12.6 39.776 13.272 ;
  LAYER M2 ;
        RECT 29.68 12.584 39.76 12.616 ;
  LAYER M2 ;
        RECT 30.284 12.584 30.356 12.616 ;
  LAYER M3 ;
        RECT 30.3 12.6 30.34 13.02 ;
  LAYER M2 ;
        RECT 30.284 13.004 30.356 13.036 ;
  LAYER M1 ;
        RECT 39.744 12.564 39.776 12.636 ;
  LAYER M2 ;
        RECT 39.724 12.584 39.796 12.616 ;
  LAYER M1 ;
        RECT 39.744 12.564 39.776 12.636 ;
  LAYER M2 ;
        RECT 39.724 12.584 39.796 12.616 ;
  LAYER M1 ;
        RECT 39.744 12.564 39.776 12.636 ;
  LAYER M2 ;
        RECT 39.724 12.584 39.796 12.616 ;
  LAYER M2 ;
        RECT 30.284 12.584 30.356 12.616 ;
  LAYER M3 ;
        RECT 30.3 12.564 30.34 12.636 ;
  LAYER M2 ;
        RECT 30.284 13.004 30.356 13.036 ;
  LAYER M3 ;
        RECT 30.3 12.984 30.34 13.056 ;
  LAYER M1 ;
        RECT 39.744 12.564 39.776 12.636 ;
  LAYER M2 ;
        RECT 39.724 12.584 39.796 12.616 ;
  LAYER M2 ;
        RECT 30.284 12.584 30.356 12.616 ;
  LAYER M3 ;
        RECT 30.3 12.564 30.34 12.636 ;
  LAYER M2 ;
        RECT 30.284 13.004 30.356 13.036 ;
  LAYER M3 ;
        RECT 30.3 12.984 30.34 13.056 ;
  LAYER M1 ;
        RECT 49.264 39.696 49.296 39.768 ;
  LAYER M2 ;
        RECT 49.244 39.716 49.316 39.748 ;
  LAYER M1 ;
        RECT 40.064 39.696 40.096 39.768 ;
  LAYER M2 ;
        RECT 40.044 39.716 40.116 39.748 ;
  LAYER M2 ;
        RECT 40.08 39.716 49.28 39.748 ;
  LAYER M2 ;
        RECT 29.484 2 29.716 2.032 ;
  LAYER M2 ;
        RECT 42.524 10.316 48.516 10.348 ;
  LAYER M2 ;
        RECT 29.884 6.872 30.116 6.904 ;
  LAYER M2 ;
        RECT 48.044 39.716 48.116 39.748 ;
  LAYER M3 ;
        RECT 48.06 39.543 48.1 39.753 ;
  LAYER M4 ;
        RECT 48.018 39.544 48.158 39.584 ;
  LAYER M5 ;
        RECT 48.064 8.484 48.128 39.564 ;
  LAYER M4 ;
        RECT 32.112 8.464 48.096 8.504 ;
  LAYER M5 ;
        RECT 32.08 4.704 32.144 8.484 ;
  LAYER M4 ;
        RECT 31.986 4.684 32.126 4.724 ;
  LAYER M3 ;
        RECT 31.98 2.016 32.02 4.704 ;
  LAYER M2 ;
        RECT 29.68 2 32 2.032 ;
  LAYER M5 ;
        RECT 48.064 10.28 48.128 10.384 ;
  LAYER M4 ;
        RECT 48.096 10.312 48.32 10.352 ;
  LAYER M3 ;
        RECT 48.3 10.227 48.34 10.437 ;
  LAYER M2 ;
        RECT 48.284 10.316 48.356 10.348 ;
  LAYER M5 ;
        RECT 32.08 6.836 32.144 6.94 ;
  LAYER M4 ;
        RECT 30.48 6.868 32.112 6.908 ;
  LAYER M3 ;
        RECT 30.46 6.783 30.5 6.993 ;
  LAYER M2 ;
        RECT 30.08 6.872 30.48 6.904 ;
  LAYER M2 ;
        RECT 31.964 2 32.036 2.032 ;
  LAYER M3 ;
        RECT 31.98 1.98 32.02 2.052 ;
  LAYER M2 ;
        RECT 48.044 39.716 48.116 39.748 ;
  LAYER M3 ;
        RECT 48.06 39.696 48.1 39.768 ;
  LAYER M3 ;
        RECT 31.98 4.664 32.02 4.744 ;
  LAYER M4 ;
        RECT 31.96 4.684 32.04 4.724 ;
  LAYER M3 ;
        RECT 48.06 39.524 48.1 39.604 ;
  LAYER M4 ;
        RECT 48.04 39.544 48.12 39.584 ;
  LAYER M4 ;
        RECT 32.072 4.684 32.152 4.724 ;
  LAYER M5 ;
        RECT 32.08 4.664 32.144 4.744 ;
  LAYER M4 ;
        RECT 32.072 8.464 32.152 8.504 ;
  LAYER M5 ;
        RECT 32.08 8.444 32.144 8.524 ;
  LAYER M4 ;
        RECT 48.056 8.464 48.136 8.504 ;
  LAYER M5 ;
        RECT 48.064 8.444 48.128 8.524 ;
  LAYER M4 ;
        RECT 48.056 39.544 48.136 39.584 ;
  LAYER M5 ;
        RECT 48.064 39.524 48.128 39.604 ;
  LAYER M2 ;
        RECT 31.964 2 32.036 2.032 ;
  LAYER M3 ;
        RECT 31.98 1.98 32.02 2.052 ;
  LAYER M4 ;
        RECT 32.072 8.464 32.152 8.504 ;
  LAYER M5 ;
        RECT 32.08 8.444 32.144 8.524 ;
  LAYER M4 ;
        RECT 48.056 8.464 48.136 8.504 ;
  LAYER M5 ;
        RECT 48.064 8.444 48.128 8.524 ;
  LAYER M2 ;
        RECT 31.964 2 32.036 2.032 ;
  LAYER M3 ;
        RECT 31.98 1.98 32.02 2.052 ;
  LAYER M2 ;
        RECT 48.284 10.316 48.356 10.348 ;
  LAYER M3 ;
        RECT 48.3 10.296 48.34 10.368 ;
  LAYER M3 ;
        RECT 48.3 10.292 48.34 10.372 ;
  LAYER M4 ;
        RECT 48.28 10.312 48.36 10.352 ;
  LAYER M4 ;
        RECT 32.072 8.464 32.152 8.504 ;
  LAYER M5 ;
        RECT 32.08 8.444 32.144 8.524 ;
  LAYER M4 ;
        RECT 48.056 8.464 48.136 8.504 ;
  LAYER M5 ;
        RECT 48.064 8.444 48.128 8.524 ;
  LAYER M4 ;
        RECT 48.056 10.312 48.136 10.352 ;
  LAYER M5 ;
        RECT 48.064 10.292 48.128 10.372 ;
  LAYER M2 ;
        RECT 31.964 2 32.036 2.032 ;
  LAYER M3 ;
        RECT 31.98 1.98 32.02 2.052 ;
  LAYER M4 ;
        RECT 32.072 8.464 32.152 8.504 ;
  LAYER M5 ;
        RECT 32.08 8.444 32.144 8.524 ;
  LAYER M4 ;
        RECT 48.056 8.464 48.136 8.504 ;
  LAYER M5 ;
        RECT 48.064 8.444 48.128 8.524 ;
  LAYER M4 ;
        RECT 48.056 10.312 48.136 10.352 ;
  LAYER M5 ;
        RECT 48.064 10.292 48.128 10.372 ;
  LAYER M2 ;
        RECT 30.444 6.872 30.516 6.904 ;
  LAYER M3 ;
        RECT 30.46 6.852 30.5 6.924 ;
  LAYER M2 ;
        RECT 31.964 2 32.036 2.032 ;
  LAYER M3 ;
        RECT 31.98 1.98 32.02 2.052 ;
  LAYER M3 ;
        RECT 30.46 6.848 30.5 6.928 ;
  LAYER M4 ;
        RECT 30.44 6.868 30.52 6.908 ;
  LAYER M4 ;
        RECT 32.072 6.868 32.152 6.908 ;
  LAYER M5 ;
        RECT 32.08 6.848 32.144 6.928 ;
  LAYER M4 ;
        RECT 32.072 8.464 32.152 8.504 ;
  LAYER M5 ;
        RECT 32.08 8.444 32.144 8.524 ;
  LAYER M4 ;
        RECT 48.056 8.464 48.136 8.504 ;
  LAYER M5 ;
        RECT 48.064 8.444 48.128 8.524 ;
  LAYER M4 ;
        RECT 48.056 10.312 48.136 10.352 ;
  LAYER M5 ;
        RECT 48.064 10.292 48.128 10.372 ;
  LAYER M2 ;
        RECT 31.964 2 32.036 2.032 ;
  LAYER M3 ;
        RECT 31.98 1.98 32.02 2.052 ;
  LAYER M4 ;
        RECT 32.072 6.868 32.152 6.908 ;
  LAYER M5 ;
        RECT 32.08 6.848 32.144 6.928 ;
  LAYER M4 ;
        RECT 32.072 8.464 32.152 8.504 ;
  LAYER M5 ;
        RECT 32.08 8.444 32.144 8.524 ;
  LAYER M4 ;
        RECT 48.056 8.464 48.136 8.504 ;
  LAYER M5 ;
        RECT 48.064 8.444 48.128 8.524 ;
  LAYER M4 ;
        RECT 48.056 10.312 48.136 10.352 ;
  LAYER M5 ;
        RECT 48.064 10.292 48.128 10.372 ;
  LAYER M1 ;
        RECT 9.584 13.236 9.616 13.308 ;
  LAYER M2 ;
        RECT 9.564 13.256 9.636 13.288 ;
  LAYER M1 ;
        RECT 18.784 13.236 18.816 13.308 ;
  LAYER M2 ;
        RECT 18.764 13.256 18.836 13.288 ;
  LAYER M2 ;
        RECT 9.6 13.256 18.8 13.288 ;
  LAYER M2 ;
        RECT 28.844 12.5 29.076 12.532 ;
  LAYER M2 ;
        RECT 28.124 13.004 28.356 13.036 ;
  LAYER M1 ;
        RECT 18.784 12.516 18.816 13.272 ;
  LAYER M2 ;
        RECT 18.8 12.5 28.88 12.532 ;
  LAYER M2 ;
        RECT 28.204 12.5 28.276 12.532 ;
  LAYER M3 ;
        RECT 28.22 12.516 28.26 13.02 ;
  LAYER M2 ;
        RECT 28.204 13.004 28.276 13.036 ;
  LAYER M1 ;
        RECT 18.784 12.48 18.816 12.552 ;
  LAYER M2 ;
        RECT 18.764 12.5 18.836 12.532 ;
  LAYER M1 ;
        RECT 18.784 12.48 18.816 12.552 ;
  LAYER M2 ;
        RECT 18.764 12.5 18.836 12.532 ;
  LAYER M1 ;
        RECT 18.784 12.48 18.816 12.552 ;
  LAYER M2 ;
        RECT 18.764 12.5 18.836 12.532 ;
  LAYER M2 ;
        RECT 28.204 12.5 28.276 12.532 ;
  LAYER M3 ;
        RECT 28.22 12.48 28.26 12.552 ;
  LAYER M2 ;
        RECT 28.204 13.004 28.276 13.036 ;
  LAYER M3 ;
        RECT 28.22 12.984 28.26 13.056 ;
  LAYER M1 ;
        RECT 18.784 12.48 18.816 12.552 ;
  LAYER M2 ;
        RECT 18.764 12.5 18.836 12.532 ;
  LAYER M2 ;
        RECT 28.204 12.5 28.276 12.532 ;
  LAYER M3 ;
        RECT 28.22 12.48 28.26 12.552 ;
  LAYER M2 ;
        RECT 28.204 13.004 28.276 13.036 ;
  LAYER M3 ;
        RECT 28.22 12.984 28.26 13.056 ;
  LAYER M1 ;
        RECT 9.264 39.696 9.296 39.768 ;
  LAYER M2 ;
        RECT 9.244 39.716 9.316 39.748 ;
  LAYER M1 ;
        RECT 18.464 39.696 18.496 39.768 ;
  LAYER M2 ;
        RECT 18.444 39.716 18.516 39.748 ;
  LAYER M2 ;
        RECT 9.28 39.716 18.48 39.748 ;
  LAYER M2 ;
        RECT 28.844 2.084 29.076 2.116 ;
  LAYER M2 ;
        RECT 10.044 10.316 16.036 10.348 ;
  LAYER M2 ;
        RECT 28.444 6.872 28.676 6.904 ;
  LAYER M2 ;
        RECT 15.964 39.716 16.036 39.748 ;
  LAYER M3 ;
        RECT 15.98 39.543 16.02 39.753 ;
  LAYER M4 ;
        RECT 15.922 39.544 16.062 39.584 ;
  LAYER M5 ;
        RECT 15.952 13.608 16.016 39.564 ;
  LAYER M4 ;
        RECT 15.922 13.588 16.062 13.628 ;
  LAYER M3 ;
        RECT 15.98 2.1 16.02 13.608 ;
  LAYER M2 ;
        RECT 16 2.084 28.88 2.116 ;
  LAYER M3 ;
        RECT 15.98 10.292 16.02 10.372 ;
  LAYER M2 ;
        RECT 15.964 10.316 16.036 10.348 ;
  LAYER M2 ;
        RECT 28.524 2.084 28.596 2.116 ;
  LAYER M3 ;
        RECT 28.54 2.1 28.58 6.888 ;
  LAYER M2 ;
        RECT 28.524 6.872 28.596 6.904 ;
  LAYER M2 ;
        RECT 15.964 2.084 16.036 2.116 ;
  LAYER M3 ;
        RECT 15.98 2.064 16.02 2.136 ;
  LAYER M2 ;
        RECT 15.964 39.716 16.036 39.748 ;
  LAYER M3 ;
        RECT 15.98 39.696 16.02 39.768 ;
  LAYER M3 ;
        RECT 15.98 13.568 16.02 13.648 ;
  LAYER M4 ;
        RECT 15.96 13.588 16.04 13.628 ;
  LAYER M3 ;
        RECT 15.98 39.524 16.02 39.604 ;
  LAYER M4 ;
        RECT 15.96 39.544 16.04 39.584 ;
  LAYER M4 ;
        RECT 15.944 13.588 16.024 13.628 ;
  LAYER M5 ;
        RECT 15.952 13.568 16.016 13.648 ;
  LAYER M4 ;
        RECT 15.944 39.544 16.024 39.584 ;
  LAYER M5 ;
        RECT 15.952 39.524 16.016 39.604 ;
  LAYER M2 ;
        RECT 15.964 2.084 16.036 2.116 ;
  LAYER M3 ;
        RECT 15.98 2.064 16.02 2.136 ;
  LAYER M2 ;
        RECT 15.964 2.084 16.036 2.116 ;
  LAYER M3 ;
        RECT 15.98 2.064 16.02 2.136 ;
  LAYER M2 ;
        RECT 15.964 10.316 16.036 10.348 ;
  LAYER M3 ;
        RECT 15.98 10.296 16.02 10.368 ;
  LAYER M2 ;
        RECT 15.964 2.084 16.036 2.116 ;
  LAYER M3 ;
        RECT 15.98 2.064 16.02 2.136 ;
  LAYER M2 ;
        RECT 15.964 10.316 16.036 10.348 ;
  LAYER M3 ;
        RECT 15.98 10.296 16.02 10.368 ;
  LAYER M2 ;
        RECT 15.964 2.084 16.036 2.116 ;
  LAYER M3 ;
        RECT 15.98 2.064 16.02 2.136 ;
  LAYER M2 ;
        RECT 15.964 10.316 16.036 10.348 ;
  LAYER M3 ;
        RECT 15.98 10.296 16.02 10.368 ;
  LAYER M2 ;
        RECT 28.524 2.084 28.596 2.116 ;
  LAYER M3 ;
        RECT 28.54 2.064 28.58 2.136 ;
  LAYER M2 ;
        RECT 28.524 6.872 28.596 6.904 ;
  LAYER M3 ;
        RECT 28.54 6.852 28.58 6.924 ;
  LAYER M2 ;
        RECT 15.964 2.084 16.036 2.116 ;
  LAYER M3 ;
        RECT 15.98 2.064 16.02 2.136 ;
  LAYER M2 ;
        RECT 15.964 10.316 16.036 10.348 ;
  LAYER M3 ;
        RECT 15.98 10.296 16.02 10.368 ;
  LAYER M2 ;
        RECT 28.524 2.084 28.596 2.116 ;
  LAYER M3 ;
        RECT 28.54 2.064 28.58 2.136 ;
  LAYER M2 ;
        RECT 28.524 6.872 28.596 6.904 ;
  LAYER M3 ;
        RECT 28.54 6.852 28.58 6.924 ;
  LAYER M2 ;
        RECT 29.324 4.856 29.556 4.888 ;
  LAYER M2 ;
        RECT 28.924 4.52 29.156 4.552 ;
  LAYER M2 ;
        RECT 42.524 4.856 48.516 4.888 ;
  LAYER M2 ;
        RECT 29.324 4.856 29.396 4.888 ;
  LAYER M3 ;
        RECT 29.34 4.536 29.38 4.872 ;
  LAYER M2 ;
        RECT 29.12 4.52 29.36 4.552 ;
  LAYER M2 ;
        RECT 29.484 4.856 29.556 4.888 ;
  LAYER M1 ;
        RECT 29.504 4.788 29.536 4.968 ;
  LAYER M2 ;
        RECT 29.52 4.772 42.56 4.804 ;
  LAYER M1 ;
        RECT 42.544 4.74 42.576 4.92 ;
  LAYER M2 ;
        RECT 42.524 4.856 42.596 4.888 ;
  LAYER M2 ;
        RECT 29.324 4.52 29.396 4.552 ;
  LAYER M3 ;
        RECT 29.34 4.5 29.38 4.572 ;
  LAYER M2 ;
        RECT 29.324 4.856 29.396 4.888 ;
  LAYER M3 ;
        RECT 29.34 4.836 29.38 4.908 ;
  LAYER M2 ;
        RECT 29.324 4.52 29.396 4.552 ;
  LAYER M3 ;
        RECT 29.34 4.5 29.38 4.572 ;
  LAYER M2 ;
        RECT 29.324 4.856 29.396 4.888 ;
  LAYER M3 ;
        RECT 29.34 4.836 29.38 4.908 ;
  LAYER M1 ;
        RECT 29.504 4.752 29.536 4.824 ;
  LAYER M2 ;
        RECT 29.484 4.772 29.556 4.804 ;
  LAYER M1 ;
        RECT 29.504 4.836 29.536 4.908 ;
  LAYER M2 ;
        RECT 29.484 4.856 29.556 4.888 ;
  LAYER M1 ;
        RECT 42.544 4.752 42.576 4.824 ;
  LAYER M2 ;
        RECT 42.524 4.772 42.596 4.804 ;
  LAYER M1 ;
        RECT 42.544 4.836 42.576 4.908 ;
  LAYER M2 ;
        RECT 42.524 4.856 42.596 4.888 ;
  LAYER M2 ;
        RECT 29.324 4.52 29.396 4.552 ;
  LAYER M3 ;
        RECT 29.34 4.5 29.38 4.572 ;
  LAYER M2 ;
        RECT 29.324 4.856 29.396 4.888 ;
  LAYER M3 ;
        RECT 29.34 4.836 29.38 4.908 ;
  LAYER M1 ;
        RECT 29.504 4.752 29.536 4.824 ;
  LAYER M2 ;
        RECT 29.484 4.772 29.556 4.804 ;
  LAYER M2 ;
        RECT 29.324 4.52 29.396 4.552 ;
  LAYER M3 ;
        RECT 29.34 4.5 29.38 4.572 ;
  LAYER M2 ;
        RECT 29.324 4.856 29.396 4.888 ;
  LAYER M3 ;
        RECT 29.34 4.836 29.38 4.908 ;
  LAYER M2 ;
        RECT 29.164 4.94 29.396 4.972 ;
  LAYER M2 ;
        RECT 29.404 4.604 29.636 4.636 ;
  LAYER M2 ;
        RECT 10.044 4.856 16.036 4.888 ;
  LAYER M2 ;
        RECT 29.36 4.94 29.44 4.972 ;
  LAYER M3 ;
        RECT 29.42 4.62 29.46 4.956 ;
  LAYER M2 ;
        RECT 29.404 4.604 29.476 4.636 ;
  LAYER M2 ;
        RECT 28.32 4.94 29.2 4.972 ;
  LAYER M3 ;
        RECT 28.3 4.851 28.34 5.061 ;
  LAYER M4 ;
        RECT 15.92 4.936 28.32 4.976 ;
  LAYER M3 ;
        RECT 15.9 4.809 15.94 5.019 ;
  LAYER M2 ;
        RECT 15.884 4.856 15.956 4.888 ;
  LAYER M2 ;
        RECT 29.404 4.604 29.476 4.636 ;
  LAYER M3 ;
        RECT 29.42 4.584 29.46 4.656 ;
  LAYER M2 ;
        RECT 29.404 4.94 29.476 4.972 ;
  LAYER M3 ;
        RECT 29.42 4.92 29.46 4.992 ;
  LAYER M2 ;
        RECT 29.404 4.604 29.476 4.636 ;
  LAYER M3 ;
        RECT 29.42 4.584 29.46 4.656 ;
  LAYER M2 ;
        RECT 29.404 4.94 29.476 4.972 ;
  LAYER M3 ;
        RECT 29.42 4.92 29.46 4.992 ;
  LAYER M2 ;
        RECT 15.884 4.856 15.956 4.888 ;
  LAYER M3 ;
        RECT 15.9 4.836 15.94 4.908 ;
  LAYER M2 ;
        RECT 28.284 4.94 28.356 4.972 ;
  LAYER M3 ;
        RECT 28.3 4.92 28.34 4.992 ;
  LAYER M2 ;
        RECT 29.404 4.604 29.476 4.636 ;
  LAYER M3 ;
        RECT 29.42 4.584 29.46 4.656 ;
  LAYER M2 ;
        RECT 29.404 4.94 29.476 4.972 ;
  LAYER M3 ;
        RECT 29.42 4.92 29.46 4.992 ;
  LAYER M3 ;
        RECT 15.9 4.916 15.94 4.996 ;
  LAYER M4 ;
        RECT 15.88 4.936 15.96 4.976 ;
  LAYER M3 ;
        RECT 28.3 4.916 28.34 4.996 ;
  LAYER M4 ;
        RECT 28.28 4.936 28.36 4.976 ;
  LAYER M2 ;
        RECT 29.404 4.604 29.476 4.636 ;
  LAYER M3 ;
        RECT 29.42 4.584 29.46 4.656 ;
  LAYER M2 ;
        RECT 29.404 4.94 29.476 4.972 ;
  LAYER M3 ;
        RECT 29.42 4.92 29.46 4.992 ;
  LAYER M2 ;
        RECT 28.844 23.588 29.716 23.62 ;
  LAYER M2 ;
        RECT 28.764 21.32 29.796 21.352 ;
  LAYER M2 ;
        RECT 29.244 23.588 29.316 23.62 ;
  LAYER M3 ;
        RECT 29.26 21.336 29.3 23.604 ;
  LAYER M2 ;
        RECT 29.244 21.32 29.316 21.352 ;
  LAYER M2 ;
        RECT 29.244 21.32 29.316 21.352 ;
  LAYER M3 ;
        RECT 29.26 21.3 29.3 21.372 ;
  LAYER M2 ;
        RECT 29.244 23.588 29.316 23.62 ;
  LAYER M3 ;
        RECT 29.26 23.568 29.3 23.64 ;
  LAYER M2 ;
        RECT 29.244 21.32 29.316 21.352 ;
  LAYER M3 ;
        RECT 29.26 21.3 29.3 21.372 ;
  LAYER M2 ;
        RECT 29.244 23.588 29.316 23.62 ;
  LAYER M3 ;
        RECT 29.26 23.568 29.3 23.64 ;
  LAYER M2 ;
        RECT 29.324 18.8 29.556 18.832 ;
  LAYER M3 ;
        RECT 29.5 16.512 29.54 18.18 ;
  LAYER M2 ;
        RECT 29.484 18.8 29.556 18.832 ;
  LAYER M3 ;
        RECT 29.5 18.144 29.54 18.816 ;
  LAYER M2 ;
        RECT 29.484 18.8 29.556 18.832 ;
  LAYER M3 ;
        RECT 29.5 18.78 29.54 18.852 ;
  LAYER M2 ;
        RECT 29.484 18.8 29.556 18.832 ;
  LAYER M3 ;
        RECT 29.5 18.78 29.54 18.852 ;
  LAYER M2 ;
        RECT 29.164 18.884 29.396 18.916 ;
  LAYER M3 ;
        RECT 29.02 16.512 29.06 18.18 ;
  LAYER M2 ;
        RECT 29.04 18.884 29.2 18.916 ;
  LAYER M3 ;
        RECT 29.02 18.144 29.06 18.9 ;
  LAYER M2 ;
        RECT 29.004 18.884 29.076 18.916 ;
  LAYER M3 ;
        RECT 29.02 18.864 29.06 18.936 ;
  LAYER M2 ;
        RECT 29.004 18.884 29.076 18.916 ;
  LAYER M3 ;
        RECT 29.02 18.864 29.06 18.936 ;
  LAYER M3 ;
        RECT 29.26 14.916 29.3 16.164 ;
  LAYER M2 ;
        RECT 29.004 21.236 29.716 21.268 ;
  LAYER M3 ;
        RECT 29.26 16.128 29.3 16.716 ;
  LAYER M2 ;
        RECT 29.22 16.7 29.42 16.732 ;
  LAYER M3 ;
        RECT 29.34 16.716 29.38 21.252 ;
  LAYER M2 ;
        RECT 29.324 21.236 29.396 21.268 ;
  LAYER M2 ;
        RECT 29.244 16.7 29.316 16.732 ;
  LAYER M3 ;
        RECT 29.26 16.68 29.3 16.752 ;
  LAYER M2 ;
        RECT 29.324 16.7 29.396 16.732 ;
  LAYER M3 ;
        RECT 29.34 16.68 29.38 16.752 ;
  LAYER M2 ;
        RECT 29.324 21.236 29.396 21.268 ;
  LAYER M3 ;
        RECT 29.34 21.216 29.38 21.288 ;
  LAYER M2 ;
        RECT 29.324 21.236 29.396 21.268 ;
  LAYER M3 ;
        RECT 29.34 21.216 29.38 21.288 ;
  LAYER M3 ;
        RECT 29.34 14.832 29.38 16.08 ;
  LAYER M2 ;
        RECT 28.844 21.152 29.556 21.184 ;
  LAYER M3 ;
        RECT 29.34 16.004 29.38 16.084 ;
  LAYER M4 ;
        RECT 29.33 16.024 29.47 16.064 ;
  LAYER M3 ;
        RECT 29.42 16.044 29.46 21.168 ;
  LAYER M2 ;
        RECT 29.404 21.152 29.476 21.184 ;
  LAYER M2 ;
        RECT 29.404 21.152 29.476 21.184 ;
  LAYER M3 ;
        RECT 29.42 21.132 29.46 21.204 ;
  LAYER M3 ;
        RECT 29.34 16.004 29.38 16.084 ;
  LAYER M4 ;
        RECT 29.32 16.024 29.4 16.064 ;
  LAYER M3 ;
        RECT 29.42 16.004 29.46 16.084 ;
  LAYER M4 ;
        RECT 29.4 16.024 29.48 16.064 ;
  LAYER M2 ;
        RECT 29.404 21.152 29.476 21.184 ;
  LAYER M3 ;
        RECT 29.42 21.132 29.46 21.204 ;
  LAYER M1 ;
        RECT 29.664 23.484 29.696 24.228 ;
  LAYER M1 ;
        RECT 29.664 24.324 29.696 24.564 ;
  LAYER M1 ;
        RECT 29.664 25.08 29.696 25.32 ;
  LAYER M1 ;
        RECT 29.744 23.484 29.776 24.228 ;
  LAYER M1 ;
        RECT 29.584 23.484 29.616 24.228 ;
  LAYER M1 ;
        RECT 29.504 23.484 29.536 24.228 ;
  LAYER M1 ;
        RECT 29.504 24.324 29.536 24.564 ;
  LAYER M1 ;
        RECT 29.504 25.08 29.536 25.32 ;
  LAYER M1 ;
        RECT 29.424 23.484 29.456 24.228 ;
  LAYER M1 ;
        RECT 29.344 23.484 29.376 24.228 ;
  LAYER M1 ;
        RECT 29.344 24.324 29.376 24.564 ;
  LAYER M1 ;
        RECT 29.344 25.08 29.376 25.32 ;
  LAYER M1 ;
        RECT 29.264 23.484 29.296 24.228 ;
  LAYER M1 ;
        RECT 29.184 23.484 29.216 24.228 ;
  LAYER M1 ;
        RECT 29.184 24.324 29.216 24.564 ;
  LAYER M1 ;
        RECT 29.184 25.08 29.216 25.32 ;
  LAYER M1 ;
        RECT 29.104 23.484 29.136 24.228 ;
  LAYER M1 ;
        RECT 29.024 23.484 29.056 24.228 ;
  LAYER M1 ;
        RECT 29.024 24.324 29.056 24.564 ;
  LAYER M1 ;
        RECT 29.024 25.08 29.056 25.32 ;
  LAYER M1 ;
        RECT 28.944 23.484 28.976 24.228 ;
  LAYER M1 ;
        RECT 28.864 23.484 28.896 24.228 ;
  LAYER M1 ;
        RECT 28.864 24.324 28.896 24.564 ;
  LAYER M1 ;
        RECT 28.864 25.08 28.896 25.32 ;
  LAYER M1 ;
        RECT 28.784 23.484 28.816 24.228 ;
  LAYER M2 ;
        RECT 29.004 23.504 29.556 23.536 ;
  LAYER M2 ;
        RECT 28.844 24.344 29.716 24.376 ;
  LAYER M2 ;
        RECT 28.844 25.184 29.716 25.216 ;
  LAYER M2 ;
        RECT 28.764 23.672 29.796 23.704 ;
  LAYER M3 ;
        RECT 29.5 23.484 29.54 24.396 ;
  LAYER M2 ;
        RECT 28.844 23.588 29.716 23.62 ;
  LAYER M3 ;
        RECT 29.34 23.652 29.38 25.236 ;
  LAYER M1 ;
        RECT 29.344 18.78 29.376 19.524 ;
  LAYER M1 ;
        RECT 29.344 19.62 29.376 19.86 ;
  LAYER M1 ;
        RECT 29.344 20.376 29.376 20.616 ;
  LAYER M1 ;
        RECT 29.424 18.78 29.456 19.524 ;
  LAYER M1 ;
        RECT 29.264 18.78 29.296 19.524 ;
  LAYER M1 ;
        RECT 29.184 18.78 29.216 19.524 ;
  LAYER M1 ;
        RECT 29.184 19.62 29.216 19.86 ;
  LAYER M1 ;
        RECT 29.184 20.376 29.216 20.616 ;
  LAYER M1 ;
        RECT 29.104 18.78 29.136 19.524 ;
  LAYER M2 ;
        RECT 29.164 20.48 29.396 20.512 ;
  LAYER M2 ;
        RECT 29.084 18.968 29.476 19 ;
  LAYER M2 ;
        RECT 29.324 18.8 29.556 18.832 ;
  LAYER M2 ;
        RECT 29.164 18.884 29.396 18.916 ;
  LAYER M2 ;
        RECT 29.164 19.64 29.396 19.672 ;
  LAYER M3 ;
        RECT 29.26 18.948 29.3 20.532 ;
  LAYER M1 ;
        RECT 29.584 16.428 29.616 17.172 ;
  LAYER M1 ;
        RECT 29.584 17.268 29.616 17.508 ;
  LAYER M1 ;
        RECT 29.584 18.024 29.616 18.264 ;
  LAYER M1 ;
        RECT 29.504 16.428 29.536 17.172 ;
  LAYER M1 ;
        RECT 29.664 16.428 29.696 17.172 ;
  LAYER M2 ;
        RECT 29.404 18.128 29.636 18.16 ;
  LAYER M2 ;
        RECT 29.484 16.532 29.716 16.564 ;
  LAYER M2 ;
        RECT 29.404 16.448 29.636 16.48 ;
  LAYER M2 ;
        RECT 29.404 17.288 29.636 17.32 ;
  LAYER M3 ;
        RECT 29.5 16.512 29.54 18.18 ;
  LAYER M1 ;
        RECT 28.944 16.428 28.976 17.172 ;
  LAYER M1 ;
        RECT 28.944 17.268 28.976 17.508 ;
  LAYER M1 ;
        RECT 28.944 18.024 28.976 18.264 ;
  LAYER M1 ;
        RECT 29.024 16.428 29.056 17.172 ;
  LAYER M1 ;
        RECT 28.864 16.428 28.896 17.172 ;
  LAYER M2 ;
        RECT 28.924 18.128 29.156 18.16 ;
  LAYER M2 ;
        RECT 28.844 16.532 29.076 16.564 ;
  LAYER M2 ;
        RECT 28.924 16.448 29.156 16.48 ;
  LAYER M2 ;
        RECT 28.924 17.288 29.156 17.32 ;
  LAYER M3 ;
        RECT 29.02 16.512 29.06 18.18 ;
  LAYER M1 ;
        RECT 28.944 15.588 28.976 16.332 ;
  LAYER M1 ;
        RECT 28.944 15.252 28.976 15.492 ;
  LAYER M1 ;
        RECT 28.944 14.412 28.976 15.156 ;
  LAYER M1 ;
        RECT 28.944 14.076 28.976 14.316 ;
  LAYER M1 ;
        RECT 28.944 13.32 28.976 13.56 ;
  LAYER M1 ;
        RECT 28.864 15.588 28.896 16.332 ;
  LAYER M1 ;
        RECT 28.864 14.412 28.896 15.156 ;
  LAYER M1 ;
        RECT 29.024 15.588 29.056 16.332 ;
  LAYER M1 ;
        RECT 29.024 14.412 29.056 15.156 ;
  LAYER M1 ;
        RECT 29.584 15.588 29.616 16.332 ;
  LAYER M1 ;
        RECT 29.584 15.252 29.616 15.492 ;
  LAYER M1 ;
        RECT 29.584 14.412 29.616 15.156 ;
  LAYER M1 ;
        RECT 29.584 14.076 29.616 14.316 ;
  LAYER M1 ;
        RECT 29.584 13.32 29.616 13.56 ;
  LAYER M1 ;
        RECT 29.504 15.588 29.536 16.332 ;
  LAYER M1 ;
        RECT 29.504 14.412 29.536 15.156 ;
  LAYER M1 ;
        RECT 29.664 15.588 29.696 16.332 ;
  LAYER M1 ;
        RECT 29.664 14.412 29.696 15.156 ;
  LAYER M2 ;
        RECT 28.924 16.28 29.156 16.312 ;
  LAYER M2 ;
        RECT 29.164 16.196 29.636 16.228 ;
  LAYER M2 ;
        RECT 28.844 16.112 29.316 16.144 ;
  LAYER M2 ;
        RECT 29.324 16.028 29.716 16.06 ;
  LAYER M2 ;
        RECT 28.924 15.44 29.636 15.472 ;
  LAYER M2 ;
        RECT 29.084 15.104 29.636 15.136 ;
  LAYER M2 ;
        RECT 28.924 15.02 29.236 15.052 ;
  LAYER M2 ;
        RECT 29.244 14.936 29.716 14.968 ;
  LAYER M2 ;
        RECT 28.844 14.852 29.396 14.884 ;
  LAYER M2 ;
        RECT 28.924 14.264 29.636 14.296 ;
  LAYER M2 ;
        RECT 28.924 13.424 29.636 13.456 ;
  LAYER M3 ;
        RECT 29.1 15.084 29.14 16.332 ;
  LAYER M3 ;
        RECT 29.18 15 29.22 16.248 ;
  LAYER M3 ;
        RECT 29.42 14.244 29.46 15.492 ;
  LAYER M3 ;
        RECT 29.26 14.916 29.3 16.164 ;
  LAYER M3 ;
        RECT 29.34 14.832 29.38 16.08 ;
  LAYER M1 ;
        RECT 28.864 21.132 28.896 21.876 ;
  LAYER M1 ;
        RECT 28.864 21.972 28.896 22.212 ;
  LAYER M1 ;
        RECT 28.864 22.728 28.896 22.968 ;
  LAYER M1 ;
        RECT 28.784 21.132 28.816 21.876 ;
  LAYER M1 ;
        RECT 28.944 21.132 28.976 21.876 ;
  LAYER M1 ;
        RECT 29.024 21.132 29.056 21.876 ;
  LAYER M1 ;
        RECT 29.024 21.972 29.056 22.212 ;
  LAYER M1 ;
        RECT 29.024 22.728 29.056 22.968 ;
  LAYER M1 ;
        RECT 29.104 21.132 29.136 21.876 ;
  LAYER M1 ;
        RECT 29.184 21.132 29.216 21.876 ;
  LAYER M1 ;
        RECT 29.184 21.972 29.216 22.212 ;
  LAYER M1 ;
        RECT 29.184 22.728 29.216 22.968 ;
  LAYER M1 ;
        RECT 29.264 21.132 29.296 21.876 ;
  LAYER M1 ;
        RECT 29.344 21.132 29.376 21.876 ;
  LAYER M1 ;
        RECT 29.344 21.972 29.376 22.212 ;
  LAYER M1 ;
        RECT 29.344 22.728 29.376 22.968 ;
  LAYER M1 ;
        RECT 29.424 21.132 29.456 21.876 ;
  LAYER M1 ;
        RECT 29.504 21.132 29.536 21.876 ;
  LAYER M1 ;
        RECT 29.504 21.972 29.536 22.212 ;
  LAYER M1 ;
        RECT 29.504 22.728 29.536 22.968 ;
  LAYER M1 ;
        RECT 29.584 21.132 29.616 21.876 ;
  LAYER M1 ;
        RECT 29.664 21.132 29.696 21.876 ;
  LAYER M1 ;
        RECT 29.664 21.972 29.696 22.212 ;
  LAYER M1 ;
        RECT 29.664 22.728 29.696 22.968 ;
  LAYER M1 ;
        RECT 29.744 21.132 29.776 21.876 ;
  LAYER M2 ;
        RECT 28.844 22.832 29.716 22.864 ;
  LAYER M2 ;
        RECT 28.844 21.152 29.556 21.184 ;
  LAYER M2 ;
        RECT 29.004 21.236 29.716 21.268 ;
  LAYER M2 ;
        RECT 28.844 21.992 29.556 22.024 ;
  LAYER M2 ;
        RECT 29.004 22.076 29.716 22.108 ;
  LAYER M2 ;
        RECT 28.764 21.32 29.796 21.352 ;
  LAYER M1 ;
        RECT 40.304 21.666 40.336 21.856 ;
  LAYER M2 ;
        RECT 40.22 21.74 40.42 21.772 ;
  LAYER M2 ;
        RECT 40.32 21.74 49.28 21.772 ;
  LAYER M1 ;
        RECT 49.264 21.72 49.296 21.792 ;
  LAYER M2 ;
        RECT 49.244 21.74 49.316 21.772 ;
  LAYER M1 ;
        RECT 49.504 30.318 49.536 30.508 ;
  LAYER M2 ;
        RECT 49.42 30.392 49.62 30.424 ;
  LAYER M1 ;
        RECT 49.504 30.408 49.536 30.576 ;
  LAYER M1 ;
        RECT 49.504 30.54 49.536 30.612 ;
  LAYER M2 ;
        RECT 49.484 30.56 49.556 30.592 ;
  LAYER M2 ;
        RECT 49.28 30.56 49.52 30.592 ;
  LAYER M1 ;
        RECT 49.264 30.54 49.296 30.612 ;
  LAYER M2 ;
        RECT 49.244 30.56 49.316 30.592 ;
  LAYER M1 ;
        RECT 49.264 39.696 49.296 39.768 ;
  LAYER M2 ;
        RECT 49.244 39.716 49.316 39.748 ;
  LAYER M1 ;
        RECT 49.264 39.396 49.296 39.732 ;
  LAYER M1 ;
        RECT 49.264 21.756 49.296 39.396 ;
  LAYER M1 ;
        RECT 31.104 30.318 31.136 30.508 ;
  LAYER M2 ;
        RECT 31.02 30.392 31.22 30.424 ;
  LAYER M2 ;
        RECT 31.12 30.392 40.08 30.424 ;
  LAYER M1 ;
        RECT 40.064 30.372 40.096 30.444 ;
  LAYER M2 ;
        RECT 40.044 30.392 40.116 30.424 ;
  LAYER M1 ;
        RECT 40.064 39.696 40.096 39.768 ;
  LAYER M2 ;
        RECT 40.044 39.716 40.116 39.748 ;
  LAYER M1 ;
        RECT 40.064 39.396 40.096 39.732 ;
  LAYER M1 ;
        RECT 40.064 30.408 40.096 39.396 ;
  LAYER M2 ;
        RECT 40.08 39.716 49.28 39.748 ;
  LAYER M1 ;
        RECT 49.504 38.97 49.536 39.16 ;
  LAYER M2 ;
        RECT 49.42 39.044 49.62 39.076 ;
  LAYER M2 ;
        RECT 49.52 39.044 58.48 39.076 ;
  LAYER M1 ;
        RECT 58.464 39.024 58.496 39.096 ;
  LAYER M2 ;
        RECT 58.444 39.044 58.516 39.076 ;
  LAYER M1 ;
        RECT 49.504 21.666 49.536 21.856 ;
  LAYER M2 ;
        RECT 49.42 21.74 49.62 21.772 ;
  LAYER M2 ;
        RECT 49.52 21.74 58.48 21.772 ;
  LAYER M1 ;
        RECT 58.464 21.72 58.496 21.792 ;
  LAYER M2 ;
        RECT 58.444 21.74 58.516 21.772 ;
  LAYER M1 ;
        RECT 58.464 39.864 58.496 39.936 ;
  LAYER M2 ;
        RECT 58.444 39.884 58.516 39.916 ;
  LAYER M1 ;
        RECT 58.464 39.396 58.496 39.9 ;
  LAYER M1 ;
        RECT 58.464 21.756 58.496 39.396 ;
  LAYER M1 ;
        RECT 31.104 21.666 31.136 21.856 ;
  LAYER M2 ;
        RECT 31.02 21.74 31.22 21.772 ;
  LAYER M1 ;
        RECT 31.104 21.756 31.136 21.924 ;
  LAYER M1 ;
        RECT 31.104 21.888 31.136 21.96 ;
  LAYER M2 ;
        RECT 31.084 21.908 31.156 21.94 ;
  LAYER M2 ;
        RECT 30.88 21.908 31.12 21.94 ;
  LAYER M1 ;
        RECT 30.864 21.888 30.896 21.96 ;
  LAYER M2 ;
        RECT 30.844 21.908 30.916 21.94 ;
  LAYER M1 ;
        RECT 31.104 38.97 31.136 39.16 ;
  LAYER M2 ;
        RECT 31.02 39.044 31.22 39.076 ;
  LAYER M1 ;
        RECT 31.104 39.06 31.136 39.228 ;
  LAYER M1 ;
        RECT 31.104 39.192 31.136 39.264 ;
  LAYER M2 ;
        RECT 31.084 39.212 31.156 39.244 ;
  LAYER M2 ;
        RECT 30.88 39.212 31.12 39.244 ;
  LAYER M1 ;
        RECT 30.864 39.192 30.896 39.264 ;
  LAYER M2 ;
        RECT 30.844 39.212 30.916 39.244 ;
  LAYER M1 ;
        RECT 30.864 39.864 30.896 39.936 ;
  LAYER M2 ;
        RECT 30.844 39.884 30.916 39.916 ;
  LAYER M1 ;
        RECT 30.864 39.396 30.896 39.9 ;
  LAYER M1 ;
        RECT 30.864 21.924 30.896 39.396 ;
  LAYER M2 ;
        RECT 30.88 39.884 58.48 39.916 ;
  LAYER M1 ;
        RECT 40.304 38.97 40.336 39.16 ;
  LAYER M2 ;
        RECT 40.22 39.044 40.42 39.076 ;
  LAYER M2 ;
        RECT 40.32 39.044 49.52 39.076 ;
  LAYER M1 ;
        RECT 49.504 38.97 49.536 39.16 ;
  LAYER M2 ;
        RECT 49.42 39.044 49.62 39.076 ;
  LAYER M1 ;
        RECT 40.304 30.318 40.336 30.508 ;
  LAYER M2 ;
        RECT 40.22 30.392 40.42 30.424 ;
  LAYER M2 ;
        RECT 40.32 30.392 49.12 30.424 ;
  LAYER M1 ;
        RECT 49.104 30.372 49.136 30.444 ;
  LAYER M2 ;
        RECT 49.084 30.392 49.156 30.424 ;
  LAYER M1 ;
        RECT 49.104 40.032 49.136 40.104 ;
  LAYER M2 ;
        RECT 49.084 40.052 49.156 40.084 ;
  LAYER M1 ;
        RECT 49.104 39.396 49.136 40.068 ;
  LAYER M1 ;
        RECT 49.104 30.408 49.136 39.396 ;
  LAYER M1 ;
        RECT 49.104 40.032 49.136 40.104 ;
  LAYER M2 ;
        RECT 49.084 40.052 49.156 40.084 ;
  LAYER M1 ;
        RECT 49.104 39.396 49.136 40.068 ;
  LAYER M1 ;
        RECT 49.104 39.06 49.136 39.396 ;
  LAYER M2 ;
        RECT 48.92 40.052 49.12 40.084 ;
  LAYER M1 ;
        RECT 48.544 13.854 48.576 14.044 ;
  LAYER M2 ;
        RECT 48.46 13.928 48.66 13.96 ;
  LAYER M2 ;
        RECT 48.56 13.928 48.96 13.96 ;
  LAYER M1 ;
        RECT 48.944 13.908 48.976 13.98 ;
  LAYER M2 ;
        RECT 48.924 13.928 48.996 13.96 ;
  LAYER M1 ;
        RECT 57.744 22.506 57.776 22.696 ;
  LAYER M2 ;
        RECT 57.66 22.58 57.86 22.612 ;
  LAYER M1 ;
        RECT 57.744 22.428 57.776 22.596 ;
  LAYER M1 ;
        RECT 57.744 22.392 57.776 22.464 ;
  LAYER M2 ;
        RECT 57.724 22.412 57.796 22.444 ;
  LAYER M2 ;
        RECT 48.96 22.412 57.76 22.444 ;
  LAYER M1 ;
        RECT 48.944 22.392 48.976 22.464 ;
  LAYER M2 ;
        RECT 48.924 22.412 48.996 22.444 ;
  LAYER M1 ;
        RECT 48.944 13.236 48.976 13.308 ;
  LAYER M2 ;
        RECT 48.924 13.256 48.996 13.288 ;
  LAYER M1 ;
        RECT 48.944 13.272 48.976 13.608 ;
  LAYER M1 ;
        RECT 48.944 13.608 48.976 22.428 ;
  LAYER M1 ;
        RECT 39.344 22.506 39.376 22.696 ;
  LAYER M2 ;
        RECT 39.26 22.58 39.46 22.612 ;
  LAYER M2 ;
        RECT 39.36 22.58 39.76 22.612 ;
  LAYER M1 ;
        RECT 39.744 22.56 39.776 22.632 ;
  LAYER M2 ;
        RECT 39.724 22.58 39.796 22.612 ;
  LAYER M1 ;
        RECT 39.744 13.236 39.776 13.308 ;
  LAYER M2 ;
        RECT 39.724 13.256 39.796 13.288 ;
  LAYER M1 ;
        RECT 39.744 13.272 39.776 13.608 ;
  LAYER M1 ;
        RECT 39.744 13.608 39.776 22.596 ;
  LAYER M2 ;
        RECT 39.76 13.256 48.96 13.288 ;
  LAYER M1 ;
        RECT 57.744 31.158 57.776 31.348 ;
  LAYER M2 ;
        RECT 57.66 31.232 57.86 31.264 ;
  LAYER M2 ;
        RECT 57.76 31.232 58.32 31.264 ;
  LAYER M1 ;
        RECT 58.304 31.212 58.336 31.284 ;
  LAYER M2 ;
        RECT 58.284 31.232 58.356 31.264 ;
  LAYER M1 ;
        RECT 57.744 13.854 57.776 14.044 ;
  LAYER M2 ;
        RECT 57.66 13.928 57.86 13.96 ;
  LAYER M2 ;
        RECT 57.76 13.928 58.32 13.96 ;
  LAYER M1 ;
        RECT 58.304 13.908 58.336 13.98 ;
  LAYER M2 ;
        RECT 58.284 13.928 58.356 13.96 ;
  LAYER M1 ;
        RECT 58.304 13.068 58.336 13.14 ;
  LAYER M2 ;
        RECT 58.284 13.088 58.356 13.12 ;
  LAYER M1 ;
        RECT 58.304 13.104 58.336 13.608 ;
  LAYER M1 ;
        RECT 58.304 13.608 58.336 31.248 ;
  LAYER M1 ;
        RECT 39.344 13.854 39.376 14.044 ;
  LAYER M2 ;
        RECT 39.26 13.928 39.46 13.96 ;
  LAYER M1 ;
        RECT 39.344 13.776 39.376 13.944 ;
  LAYER M1 ;
        RECT 39.344 13.74 39.376 13.812 ;
  LAYER M2 ;
        RECT 39.324 13.76 39.396 13.792 ;
  LAYER M2 ;
        RECT 30.72 13.76 39.36 13.792 ;
  LAYER M1 ;
        RECT 30.704 13.74 30.736 13.812 ;
  LAYER M2 ;
        RECT 30.684 13.76 30.756 13.792 ;
  LAYER M1 ;
        RECT 39.344 31.158 39.376 31.348 ;
  LAYER M2 ;
        RECT 39.26 31.232 39.46 31.264 ;
  LAYER M1 ;
        RECT 39.344 31.08 39.376 31.248 ;
  LAYER M1 ;
        RECT 39.344 31.044 39.376 31.116 ;
  LAYER M2 ;
        RECT 39.324 31.064 39.396 31.096 ;
  LAYER M2 ;
        RECT 30.72 31.064 39.36 31.096 ;
  LAYER M1 ;
        RECT 30.704 31.044 30.736 31.116 ;
  LAYER M2 ;
        RECT 30.684 31.064 30.756 31.096 ;
  LAYER M1 ;
        RECT 30.704 13.068 30.736 13.14 ;
  LAYER M2 ;
        RECT 30.684 13.088 30.756 13.12 ;
  LAYER M1 ;
        RECT 30.704 13.104 30.736 13.608 ;
  LAYER M1 ;
        RECT 30.704 13.608 30.736 31.08 ;
  LAYER M2 ;
        RECT 30.72 13.088 58.32 13.12 ;
  LAYER M1 ;
        RECT 48.544 31.158 48.576 31.348 ;
  LAYER M2 ;
        RECT 48.46 31.232 48.66 31.264 ;
  LAYER M2 ;
        RECT 48.56 31.232 57.76 31.264 ;
  LAYER M1 ;
        RECT 57.744 31.158 57.776 31.348 ;
  LAYER M2 ;
        RECT 57.66 31.232 57.86 31.264 ;
  LAYER M1 ;
        RECT 48.544 22.506 48.576 22.696 ;
  LAYER M2 ;
        RECT 48.46 22.58 48.66 22.612 ;
  LAYER M2 ;
        RECT 48.56 22.58 48.8 22.612 ;
  LAYER M1 ;
        RECT 48.784 22.56 48.816 22.632 ;
  LAYER M2 ;
        RECT 48.764 22.58 48.836 22.612 ;
  LAYER M1 ;
        RECT 48.784 12.9 48.816 12.972 ;
  LAYER M2 ;
        RECT 48.764 12.92 48.836 12.952 ;
  LAYER M1 ;
        RECT 48.784 12.936 48.816 13.608 ;
  LAYER M1 ;
        RECT 48.784 13.608 48.816 22.596 ;
  LAYER M1 ;
        RECT 48.784 12.9 48.816 12.972 ;
  LAYER M2 ;
        RECT 48.764 12.92 48.836 12.952 ;
  LAYER M1 ;
        RECT 48.784 12.936 48.816 13.608 ;
  LAYER M1 ;
        RECT 48.784 13.608 48.816 31.248 ;
  LAYER M2 ;
        RECT 48.6 12.92 48.8 12.952 ;
  LAYER M1 ;
        RECT 49.44 31.08 57.84 39.228 ;
  LAYER M2 ;
        RECT 49.44 31.08 57.84 39.228 ;
  LAYER M3 ;
        RECT 49.44 31.08 57.84 39.228 ;
  LAYER M1 ;
        RECT 49.44 22.428 57.84 30.576 ;
  LAYER M2 ;
        RECT 49.44 22.428 57.84 30.576 ;
  LAYER M3 ;
        RECT 49.44 22.428 57.84 30.576 ;
  LAYER M1 ;
        RECT 49.44 13.776 57.84 21.924 ;
  LAYER M2 ;
        RECT 49.44 13.776 57.84 21.924 ;
  LAYER M3 ;
        RECT 49.44 13.776 57.84 21.924 ;
  LAYER M1 ;
        RECT 40.24 31.08 48.64 39.228 ;
  LAYER M2 ;
        RECT 40.24 31.08 48.64 39.228 ;
  LAYER M3 ;
        RECT 40.24 31.08 48.64 39.228 ;
  LAYER M1 ;
        RECT 40.24 22.428 48.64 30.576 ;
  LAYER M2 ;
        RECT 40.24 22.428 48.64 30.576 ;
  LAYER M3 ;
        RECT 40.24 22.428 48.64 30.576 ;
  LAYER M1 ;
        RECT 40.24 13.776 48.64 21.924 ;
  LAYER M2 ;
        RECT 40.24 13.776 48.64 21.924 ;
  LAYER M3 ;
        RECT 40.24 13.776 48.64 21.924 ;
  LAYER M1 ;
        RECT 31.04 31.08 39.44 39.228 ;
  LAYER M2 ;
        RECT 31.04 31.08 39.44 39.228 ;
  LAYER M3 ;
        RECT 31.04 31.08 39.44 39.228 ;
  LAYER M1 ;
        RECT 31.04 22.428 39.44 30.576 ;
  LAYER M2 ;
        RECT 31.04 22.428 39.44 30.576 ;
  LAYER M3 ;
        RECT 31.04 22.428 39.44 30.576 ;
  LAYER M1 ;
        RECT 31.04 13.776 39.44 21.924 ;
  LAYER M2 ;
        RECT 31.04 13.776 39.44 21.924 ;
  LAYER M3 ;
        RECT 31.04 13.776 39.44 21.924 ;
  LAYER M1 ;
        RECT 48.944 13.236 48.976 13.308 ;
  LAYER M2 ;
        RECT 48.924 13.256 48.996 13.288 ;
  LAYER M1 ;
        RECT 39.744 13.236 39.776 13.308 ;
  LAYER M2 ;
        RECT 39.724 13.256 39.796 13.288 ;
  LAYER M2 ;
        RECT 39.76 13.256 48.96 13.288 ;
  LAYER M1 ;
        RECT 58.304 13.068 58.336 13.14 ;
  LAYER M2 ;
        RECT 58.284 13.088 58.356 13.12 ;
  LAYER M1 ;
        RECT 30.704 13.068 30.736 13.14 ;
  LAYER M2 ;
        RECT 30.684 13.088 30.756 13.12 ;
  LAYER M2 ;
        RECT 30.72 13.088 58.32 13.12 ;
  LAYER M1 ;
        RECT 49.264 39.696 49.296 39.768 ;
  LAYER M2 ;
        RECT 49.244 39.716 49.316 39.748 ;
  LAYER M1 ;
        RECT 40.064 39.696 40.096 39.768 ;
  LAYER M2 ;
        RECT 40.044 39.716 40.116 39.748 ;
  LAYER M2 ;
        RECT 40.08 39.716 49.28 39.748 ;
  LAYER M1 ;
        RECT 58.464 39.864 58.496 39.936 ;
  LAYER M2 ;
        RECT 58.444 39.884 58.516 39.916 ;
  LAYER M1 ;
        RECT 30.864 39.864 30.896 39.936 ;
  LAYER M2 ;
        RECT 30.844 39.884 30.916 39.916 ;
  LAYER M2 ;
        RECT 30.88 39.884 58.48 39.916 ;
  LAYER M1 ;
        RECT 18.224 21.666 18.256 21.856 ;
  LAYER M2 ;
        RECT 18.14 21.74 18.34 21.772 ;
  LAYER M2 ;
        RECT 9.28 21.74 18.24 21.772 ;
  LAYER M1 ;
        RECT 9.264 21.72 9.296 21.792 ;
  LAYER M2 ;
        RECT 9.244 21.74 9.316 21.772 ;
  LAYER M1 ;
        RECT 9.024 30.318 9.056 30.508 ;
  LAYER M2 ;
        RECT 8.94 30.392 9.14 30.424 ;
  LAYER M1 ;
        RECT 9.024 30.408 9.056 30.576 ;
  LAYER M1 ;
        RECT 9.024 30.54 9.056 30.612 ;
  LAYER M2 ;
        RECT 9.004 30.56 9.076 30.592 ;
  LAYER M2 ;
        RECT 9.04 30.56 9.28 30.592 ;
  LAYER M1 ;
        RECT 9.264 30.54 9.296 30.612 ;
  LAYER M2 ;
        RECT 9.244 30.56 9.316 30.592 ;
  LAYER M1 ;
        RECT 9.264 39.696 9.296 39.768 ;
  LAYER M2 ;
        RECT 9.244 39.716 9.316 39.748 ;
  LAYER M1 ;
        RECT 9.264 39.396 9.296 39.732 ;
  LAYER M1 ;
        RECT 9.264 21.756 9.296 39.396 ;
  LAYER M1 ;
        RECT 27.424 30.318 27.456 30.508 ;
  LAYER M2 ;
        RECT 27.34 30.392 27.54 30.424 ;
  LAYER M2 ;
        RECT 18.48 30.392 27.44 30.424 ;
  LAYER M1 ;
        RECT 18.464 30.372 18.496 30.444 ;
  LAYER M2 ;
        RECT 18.444 30.392 18.516 30.424 ;
  LAYER M1 ;
        RECT 18.464 39.696 18.496 39.768 ;
  LAYER M2 ;
        RECT 18.444 39.716 18.516 39.748 ;
  LAYER M1 ;
        RECT 18.464 39.396 18.496 39.732 ;
  LAYER M1 ;
        RECT 18.464 30.408 18.496 39.396 ;
  LAYER M2 ;
        RECT 9.28 39.716 18.48 39.748 ;
  LAYER M1 ;
        RECT 9.024 38.97 9.056 39.16 ;
  LAYER M2 ;
        RECT 8.94 39.044 9.14 39.076 ;
  LAYER M2 ;
        RECT 0.08 39.044 9.04 39.076 ;
  LAYER M1 ;
        RECT 0.064 39.024 0.096 39.096 ;
  LAYER M2 ;
        RECT 0.044 39.044 0.116 39.076 ;
  LAYER M1 ;
        RECT 9.024 21.666 9.056 21.856 ;
  LAYER M2 ;
        RECT 8.94 21.74 9.14 21.772 ;
  LAYER M2 ;
        RECT 0.08 21.74 9.04 21.772 ;
  LAYER M1 ;
        RECT 0.064 21.72 0.096 21.792 ;
  LAYER M2 ;
        RECT 0.044 21.74 0.116 21.772 ;
  LAYER M1 ;
        RECT 0.064 39.864 0.096 39.936 ;
  LAYER M2 ;
        RECT 0.044 39.884 0.116 39.916 ;
  LAYER M1 ;
        RECT 0.064 39.396 0.096 39.9 ;
  LAYER M1 ;
        RECT 0.064 21.756 0.096 39.396 ;
  LAYER M1 ;
        RECT 27.424 21.666 27.456 21.856 ;
  LAYER M2 ;
        RECT 27.34 21.74 27.54 21.772 ;
  LAYER M1 ;
        RECT 27.424 21.756 27.456 21.924 ;
  LAYER M1 ;
        RECT 27.424 21.888 27.456 21.96 ;
  LAYER M2 ;
        RECT 27.404 21.908 27.476 21.94 ;
  LAYER M2 ;
        RECT 27.44 21.908 27.68 21.94 ;
  LAYER M1 ;
        RECT 27.664 21.888 27.696 21.96 ;
  LAYER M2 ;
        RECT 27.644 21.908 27.716 21.94 ;
  LAYER M1 ;
        RECT 27.424 38.97 27.456 39.16 ;
  LAYER M2 ;
        RECT 27.34 39.044 27.54 39.076 ;
  LAYER M1 ;
        RECT 27.424 39.06 27.456 39.228 ;
  LAYER M1 ;
        RECT 27.424 39.192 27.456 39.264 ;
  LAYER M2 ;
        RECT 27.404 39.212 27.476 39.244 ;
  LAYER M2 ;
        RECT 27.44 39.212 27.68 39.244 ;
  LAYER M1 ;
        RECT 27.664 39.192 27.696 39.264 ;
  LAYER M2 ;
        RECT 27.644 39.212 27.716 39.244 ;
  LAYER M1 ;
        RECT 27.664 39.864 27.696 39.936 ;
  LAYER M2 ;
        RECT 27.644 39.884 27.716 39.916 ;
  LAYER M1 ;
        RECT 27.664 39.396 27.696 39.9 ;
  LAYER M1 ;
        RECT 27.664 21.924 27.696 39.396 ;
  LAYER M2 ;
        RECT 0.08 39.884 27.68 39.916 ;
  LAYER M1 ;
        RECT 18.224 38.97 18.256 39.16 ;
  LAYER M2 ;
        RECT 18.14 39.044 18.34 39.076 ;
  LAYER M2 ;
        RECT 9.04 39.044 18.24 39.076 ;
  LAYER M1 ;
        RECT 9.024 38.97 9.056 39.16 ;
  LAYER M2 ;
        RECT 8.94 39.044 9.14 39.076 ;
  LAYER M1 ;
        RECT 18.224 30.318 18.256 30.508 ;
  LAYER M2 ;
        RECT 18.14 30.392 18.34 30.424 ;
  LAYER M2 ;
        RECT 9.44 30.392 18.24 30.424 ;
  LAYER M1 ;
        RECT 9.424 30.372 9.456 30.444 ;
  LAYER M2 ;
        RECT 9.404 30.392 9.476 30.424 ;
  LAYER M1 ;
        RECT 9.424 40.032 9.456 40.104 ;
  LAYER M2 ;
        RECT 9.404 40.052 9.476 40.084 ;
  LAYER M1 ;
        RECT 9.424 39.396 9.456 40.068 ;
  LAYER M1 ;
        RECT 9.424 30.408 9.456 39.396 ;
  LAYER M1 ;
        RECT 9.424 40.032 9.456 40.104 ;
  LAYER M2 ;
        RECT 9.404 40.052 9.476 40.084 ;
  LAYER M1 ;
        RECT 9.424 39.396 9.456 40.068 ;
  LAYER M1 ;
        RECT 9.424 39.06 9.456 39.396 ;
  LAYER M2 ;
        RECT 9.44 40.052 9.64 40.084 ;
  LAYER M1 ;
        RECT 9.984 13.854 10.016 14.044 ;
  LAYER M2 ;
        RECT 9.9 13.928 10.1 13.96 ;
  LAYER M2 ;
        RECT 9.6 13.928 10 13.96 ;
  LAYER M1 ;
        RECT 9.584 13.908 9.616 13.98 ;
  LAYER M2 ;
        RECT 9.564 13.928 9.636 13.96 ;
  LAYER M1 ;
        RECT 0.784 22.506 0.816 22.696 ;
  LAYER M2 ;
        RECT 0.7 22.58 0.9 22.612 ;
  LAYER M1 ;
        RECT 0.784 22.428 0.816 22.596 ;
  LAYER M1 ;
        RECT 0.784 22.392 0.816 22.464 ;
  LAYER M2 ;
        RECT 0.764 22.412 0.836 22.444 ;
  LAYER M2 ;
        RECT 0.8 22.412 9.6 22.444 ;
  LAYER M1 ;
        RECT 9.584 22.392 9.616 22.464 ;
  LAYER M2 ;
        RECT 9.564 22.412 9.636 22.444 ;
  LAYER M1 ;
        RECT 9.584 13.236 9.616 13.308 ;
  LAYER M2 ;
        RECT 9.564 13.256 9.636 13.288 ;
  LAYER M1 ;
        RECT 9.584 13.272 9.616 13.608 ;
  LAYER M1 ;
        RECT 9.584 13.608 9.616 22.428 ;
  LAYER M1 ;
        RECT 19.184 22.506 19.216 22.696 ;
  LAYER M2 ;
        RECT 19.1 22.58 19.3 22.612 ;
  LAYER M2 ;
        RECT 18.8 22.58 19.2 22.612 ;
  LAYER M1 ;
        RECT 18.784 22.56 18.816 22.632 ;
  LAYER M2 ;
        RECT 18.764 22.58 18.836 22.612 ;
  LAYER M1 ;
        RECT 18.784 13.236 18.816 13.308 ;
  LAYER M2 ;
        RECT 18.764 13.256 18.836 13.288 ;
  LAYER M1 ;
        RECT 18.784 13.272 18.816 13.608 ;
  LAYER M1 ;
        RECT 18.784 13.608 18.816 22.596 ;
  LAYER M2 ;
        RECT 9.6 13.256 18.8 13.288 ;
  LAYER M1 ;
        RECT 0.784 31.158 0.816 31.348 ;
  LAYER M2 ;
        RECT 0.7 31.232 0.9 31.264 ;
  LAYER M2 ;
        RECT 0.24 31.232 0.8 31.264 ;
  LAYER M1 ;
        RECT 0.224 31.212 0.256 31.284 ;
  LAYER M2 ;
        RECT 0.204 31.232 0.276 31.264 ;
  LAYER M1 ;
        RECT 0.784 13.854 0.816 14.044 ;
  LAYER M2 ;
        RECT 0.7 13.928 0.9 13.96 ;
  LAYER M2 ;
        RECT 0.24 13.928 0.8 13.96 ;
  LAYER M1 ;
        RECT 0.224 13.908 0.256 13.98 ;
  LAYER M2 ;
        RECT 0.204 13.928 0.276 13.96 ;
  LAYER M1 ;
        RECT 0.224 13.068 0.256 13.14 ;
  LAYER M2 ;
        RECT 0.204 13.088 0.276 13.12 ;
  LAYER M1 ;
        RECT 0.224 13.104 0.256 13.608 ;
  LAYER M1 ;
        RECT 0.224 13.608 0.256 31.248 ;
  LAYER M1 ;
        RECT 19.184 13.854 19.216 14.044 ;
  LAYER M2 ;
        RECT 19.1 13.928 19.3 13.96 ;
  LAYER M1 ;
        RECT 19.184 13.776 19.216 13.944 ;
  LAYER M1 ;
        RECT 19.184 13.74 19.216 13.812 ;
  LAYER M2 ;
        RECT 19.164 13.76 19.236 13.792 ;
  LAYER M2 ;
        RECT 19.2 13.76 27.84 13.792 ;
  LAYER M1 ;
        RECT 27.824 13.74 27.856 13.812 ;
  LAYER M2 ;
        RECT 27.804 13.76 27.876 13.792 ;
  LAYER M1 ;
        RECT 19.184 31.158 19.216 31.348 ;
  LAYER M2 ;
        RECT 19.1 31.232 19.3 31.264 ;
  LAYER M1 ;
        RECT 19.184 31.08 19.216 31.248 ;
  LAYER M1 ;
        RECT 19.184 31.044 19.216 31.116 ;
  LAYER M2 ;
        RECT 19.164 31.064 19.236 31.096 ;
  LAYER M2 ;
        RECT 19.2 31.064 27.84 31.096 ;
  LAYER M1 ;
        RECT 27.824 31.044 27.856 31.116 ;
  LAYER M2 ;
        RECT 27.804 31.064 27.876 31.096 ;
  LAYER M1 ;
        RECT 27.824 13.068 27.856 13.14 ;
  LAYER M2 ;
        RECT 27.804 13.088 27.876 13.12 ;
  LAYER M1 ;
        RECT 27.824 13.104 27.856 13.608 ;
  LAYER M1 ;
        RECT 27.824 13.608 27.856 31.08 ;
  LAYER M2 ;
        RECT 0.24 13.088 27.84 13.12 ;
  LAYER M1 ;
        RECT 9.984 31.158 10.016 31.348 ;
  LAYER M2 ;
        RECT 9.9 31.232 10.1 31.264 ;
  LAYER M2 ;
        RECT 0.8 31.232 10 31.264 ;
  LAYER M1 ;
        RECT 0.784 31.158 0.816 31.348 ;
  LAYER M2 ;
        RECT 0.7 31.232 0.9 31.264 ;
  LAYER M1 ;
        RECT 9.984 22.506 10.016 22.696 ;
  LAYER M2 ;
        RECT 9.9 22.58 10.1 22.612 ;
  LAYER M2 ;
        RECT 9.76 22.58 10 22.612 ;
  LAYER M1 ;
        RECT 9.744 22.56 9.776 22.632 ;
  LAYER M2 ;
        RECT 9.724 22.58 9.796 22.612 ;
  LAYER M1 ;
        RECT 9.744 12.9 9.776 12.972 ;
  LAYER M2 ;
        RECT 9.724 12.92 9.796 12.952 ;
  LAYER M1 ;
        RECT 9.744 12.936 9.776 13.608 ;
  LAYER M1 ;
        RECT 9.744 13.608 9.776 22.596 ;
  LAYER M1 ;
        RECT 9.744 12.9 9.776 12.972 ;
  LAYER M2 ;
        RECT 9.724 12.92 9.796 12.952 ;
  LAYER M1 ;
        RECT 9.744 12.936 9.776 13.608 ;
  LAYER M1 ;
        RECT 9.744 13.608 9.776 31.248 ;
  LAYER M2 ;
        RECT 9.76 12.92 9.96 12.952 ;
  LAYER M1 ;
        RECT 0.72 31.08 9.12 39.228 ;
  LAYER M2 ;
        RECT 0.72 31.08 9.12 39.228 ;
  LAYER M3 ;
        RECT 0.72 31.08 9.12 39.228 ;
  LAYER M1 ;
        RECT 0.72 22.428 9.12 30.576 ;
  LAYER M2 ;
        RECT 0.72 22.428 9.12 30.576 ;
  LAYER M3 ;
        RECT 0.72 22.428 9.12 30.576 ;
  LAYER M1 ;
        RECT 0.72 13.776 9.12 21.924 ;
  LAYER M2 ;
        RECT 0.72 13.776 9.12 21.924 ;
  LAYER M3 ;
        RECT 0.72 13.776 9.12 21.924 ;
  LAYER M1 ;
        RECT 9.92 31.08 18.32 39.228 ;
  LAYER M2 ;
        RECT 9.92 31.08 18.32 39.228 ;
  LAYER M3 ;
        RECT 9.92 31.08 18.32 39.228 ;
  LAYER M1 ;
        RECT 9.92 22.428 18.32 30.576 ;
  LAYER M2 ;
        RECT 9.92 22.428 18.32 30.576 ;
  LAYER M3 ;
        RECT 9.92 22.428 18.32 30.576 ;
  LAYER M1 ;
        RECT 9.92 13.776 18.32 21.924 ;
  LAYER M2 ;
        RECT 9.92 13.776 18.32 21.924 ;
  LAYER M3 ;
        RECT 9.92 13.776 18.32 21.924 ;
  LAYER M1 ;
        RECT 19.12 31.08 27.52 39.228 ;
  LAYER M2 ;
        RECT 19.12 31.08 27.52 39.228 ;
  LAYER M3 ;
        RECT 19.12 31.08 27.52 39.228 ;
  LAYER M1 ;
        RECT 19.12 22.428 27.52 30.576 ;
  LAYER M2 ;
        RECT 19.12 22.428 27.52 30.576 ;
  LAYER M3 ;
        RECT 19.12 22.428 27.52 30.576 ;
  LAYER M1 ;
        RECT 19.12 13.776 27.52 21.924 ;
  LAYER M2 ;
        RECT 19.12 13.776 27.52 21.924 ;
  LAYER M3 ;
        RECT 19.12 13.776 27.52 21.924 ;
  LAYER M1 ;
        RECT 9.584 13.236 9.616 13.308 ;
  LAYER M2 ;
        RECT 9.564 13.256 9.636 13.288 ;
  LAYER M1 ;
        RECT 18.784 13.236 18.816 13.308 ;
  LAYER M2 ;
        RECT 18.764 13.256 18.836 13.288 ;
  LAYER M2 ;
        RECT 9.6 13.256 18.8 13.288 ;
  LAYER M1 ;
        RECT 0.224 13.068 0.256 13.14 ;
  LAYER M2 ;
        RECT 0.204 13.088 0.276 13.12 ;
  LAYER M1 ;
        RECT 27.824 13.068 27.856 13.14 ;
  LAYER M2 ;
        RECT 27.804 13.088 27.876 13.12 ;
  LAYER M2 ;
        RECT 0.24 13.088 27.84 13.12 ;
  LAYER M1 ;
        RECT 9.264 39.696 9.296 39.768 ;
  LAYER M2 ;
        RECT 9.244 39.716 9.316 39.748 ;
  LAYER M1 ;
        RECT 18.464 39.696 18.496 39.768 ;
  LAYER M2 ;
        RECT 18.444 39.716 18.516 39.748 ;
  LAYER M2 ;
        RECT 9.28 39.716 18.48 39.748 ;
  LAYER M1 ;
        RECT 0.064 39.864 0.096 39.936 ;
  LAYER M2 ;
        RECT 0.044 39.884 0.116 39.916 ;
  LAYER M1 ;
        RECT 27.664 39.864 27.696 39.936 ;
  LAYER M2 ;
        RECT 27.644 39.884 27.716 39.916 ;
  LAYER M2 ;
        RECT 0.08 39.884 27.68 39.916 ;
  LAYER M1 ;
        RECT 29.344 4.836 29.376 5.58 ;
  LAYER M1 ;
        RECT 29.344 5.676 29.376 5.916 ;
  LAYER M1 ;
        RECT 29.344 6.432 29.376 6.672 ;
  LAYER M1 ;
        RECT 29.424 4.836 29.456 5.58 ;
  LAYER M1 ;
        RECT 29.264 4.836 29.296 5.58 ;
  LAYER M1 ;
        RECT 29.184 4.836 29.216 5.58 ;
  LAYER M1 ;
        RECT 29.184 5.676 29.216 5.916 ;
  LAYER M1 ;
        RECT 29.184 6.432 29.216 6.672 ;
  LAYER M1 ;
        RECT 29.104 4.836 29.136 5.58 ;
  LAYER M2 ;
        RECT 29.164 6.536 29.396 6.568 ;
  LAYER M2 ;
        RECT 29.324 4.856 29.556 4.888 ;
  LAYER M2 ;
        RECT 29.164 4.94 29.396 4.972 ;
  LAYER M2 ;
        RECT 29.164 5.696 29.396 5.728 ;
  LAYER M2 ;
        RECT 29.084 5.024 29.476 5.056 ;
  LAYER M1 ;
        RECT 29.584 12.06 29.616 12.804 ;
  LAYER M1 ;
        RECT 29.584 11.724 29.616 11.964 ;
  LAYER M1 ;
        RECT 29.584 10.968 29.616 11.208 ;
  LAYER M1 ;
        RECT 29.664 12.06 29.696 12.804 ;
  LAYER M1 ;
        RECT 29.504 12.06 29.536 12.804 ;
  LAYER M1 ;
        RECT 28.944 12.06 28.976 12.804 ;
  LAYER M1 ;
        RECT 28.944 11.724 28.976 11.964 ;
  LAYER M1 ;
        RECT 28.944 10.968 28.976 11.208 ;
  LAYER M1 ;
        RECT 29.024 12.06 29.056 12.804 ;
  LAYER M1 ;
        RECT 28.864 12.06 28.896 12.804 ;
  LAYER M2 ;
        RECT 28.924 11.072 29.636 11.104 ;
  LAYER M2 ;
        RECT 29.404 12.752 29.636 12.784 ;
  LAYER M2 ;
        RECT 28.924 12.668 29.156 12.7 ;
  LAYER M2 ;
        RECT 28.924 11.912 29.636 11.944 ;
  LAYER M2 ;
        RECT 29.484 12.584 29.716 12.616 ;
  LAYER M2 ;
        RECT 28.844 12.5 29.076 12.532 ;
  LAYER M1 ;
        RECT 28.944 1.56 28.976 2.304 ;
  LAYER M1 ;
        RECT 28.944 1.224 28.976 1.464 ;
  LAYER M1 ;
        RECT 28.944 0.468 28.976 0.708 ;
  LAYER M1 ;
        RECT 28.864 1.56 28.896 2.304 ;
  LAYER M1 ;
        RECT 29.024 1.56 29.056 2.304 ;
  LAYER M1 ;
        RECT 29.584 1.56 29.616 2.304 ;
  LAYER M1 ;
        RECT 29.584 1.224 29.616 1.464 ;
  LAYER M1 ;
        RECT 29.584 0.468 29.616 0.708 ;
  LAYER M1 ;
        RECT 29.504 1.56 29.536 2.304 ;
  LAYER M1 ;
        RECT 29.664 1.56 29.696 2.304 ;
  LAYER M2 ;
        RECT 28.924 0.572 29.636 0.604 ;
  LAYER M2 ;
        RECT 28.924 2.252 29.156 2.284 ;
  LAYER M2 ;
        RECT 29.404 2.168 29.636 2.2 ;
  LAYER M2 ;
        RECT 28.924 1.412 29.636 1.444 ;
  LAYER M2 ;
        RECT 28.844 2.084 29.076 2.116 ;
  LAYER M2 ;
        RECT 29.484 2 29.716 2.032 ;
  LAYER M1 ;
        RECT 29.584 3.912 29.616 4.656 ;
  LAYER M1 ;
        RECT 29.584 3.576 29.616 3.816 ;
  LAYER M1 ;
        RECT 29.584 2.82 29.616 3.06 ;
  LAYER M1 ;
        RECT 29.664 3.912 29.696 4.656 ;
  LAYER M1 ;
        RECT 29.504 3.912 29.536 4.656 ;
  LAYER M1 ;
        RECT 28.944 3.912 28.976 4.656 ;
  LAYER M1 ;
        RECT 28.944 3.576 28.976 3.816 ;
  LAYER M1 ;
        RECT 28.944 2.82 28.976 3.06 ;
  LAYER M1 ;
        RECT 29.024 3.912 29.056 4.656 ;
  LAYER M1 ;
        RECT 28.864 3.912 28.896 4.656 ;
  LAYER M2 ;
        RECT 28.924 2.924 29.636 2.956 ;
  LAYER M2 ;
        RECT 29.404 4.604 29.636 4.636 ;
  LAYER M2 ;
        RECT 28.924 4.52 29.156 4.552 ;
  LAYER M2 ;
        RECT 28.924 3.764 29.636 3.796 ;
  LAYER M2 ;
        RECT 29.484 4.436 29.716 4.468 ;
  LAYER M2 ;
        RECT 28.844 4.352 29.076 4.384 ;
  LAYER M1 ;
        RECT 42.784 4.836 42.816 10.368 ;
  LAYER M1 ;
        RECT 42.848 4.836 42.88 10.368 ;
  LAYER M1 ;
        RECT 42.912 4.836 42.944 10.368 ;
  LAYER M1 ;
        RECT 42.976 4.836 43.008 10.368 ;
  LAYER M1 ;
        RECT 43.04 4.836 43.072 10.368 ;
  LAYER M1 ;
        RECT 43.104 4.836 43.136 10.368 ;
  LAYER M1 ;
        RECT 43.168 4.836 43.2 10.368 ;
  LAYER M1 ;
        RECT 43.232 4.836 43.264 10.368 ;
  LAYER M1 ;
        RECT 43.296 4.836 43.328 10.368 ;
  LAYER M1 ;
        RECT 43.36 4.836 43.392 10.368 ;
  LAYER M1 ;
        RECT 43.424 4.836 43.456 10.368 ;
  LAYER M1 ;
        RECT 43.488 4.836 43.52 10.368 ;
  LAYER M1 ;
        RECT 43.552 4.836 43.584 10.368 ;
  LAYER M1 ;
        RECT 43.616 4.836 43.648 10.368 ;
  LAYER M1 ;
        RECT 43.68 4.836 43.712 10.368 ;
  LAYER M1 ;
        RECT 43.744 4.836 43.776 10.368 ;
  LAYER M1 ;
        RECT 43.808 4.836 43.84 10.368 ;
  LAYER M1 ;
        RECT 43.872 4.836 43.904 10.368 ;
  LAYER M1 ;
        RECT 43.936 4.836 43.968 10.368 ;
  LAYER M1 ;
        RECT 44 4.836 44.032 10.368 ;
  LAYER M1 ;
        RECT 44.064 4.836 44.096 10.368 ;
  LAYER M1 ;
        RECT 44.128 4.836 44.16 10.368 ;
  LAYER M1 ;
        RECT 44.192 4.836 44.224 10.368 ;
  LAYER M1 ;
        RECT 44.256 4.836 44.288 10.368 ;
  LAYER M1 ;
        RECT 44.32 4.836 44.352 10.368 ;
  LAYER M1 ;
        RECT 44.384 4.836 44.416 10.368 ;
  LAYER M1 ;
        RECT 44.448 4.836 44.48 10.368 ;
  LAYER M1 ;
        RECT 44.512 4.836 44.544 10.368 ;
  LAYER M1 ;
        RECT 44.576 4.836 44.608 10.368 ;
  LAYER M1 ;
        RECT 44.64 4.836 44.672 10.368 ;
  LAYER M1 ;
        RECT 44.704 4.836 44.736 10.368 ;
  LAYER M1 ;
        RECT 44.768 4.836 44.8 10.368 ;
  LAYER M1 ;
        RECT 44.832 4.836 44.864 10.368 ;
  LAYER M1 ;
        RECT 44.896 4.836 44.928 10.368 ;
  LAYER M1 ;
        RECT 44.96 4.836 44.992 10.368 ;
  LAYER M1 ;
        RECT 45.024 4.836 45.056 10.368 ;
  LAYER M1 ;
        RECT 45.088 4.836 45.12 10.368 ;
  LAYER M1 ;
        RECT 45.152 4.836 45.184 10.368 ;
  LAYER M1 ;
        RECT 45.216 4.836 45.248 10.368 ;
  LAYER M1 ;
        RECT 45.28 4.836 45.312 10.368 ;
  LAYER M1 ;
        RECT 45.344 4.836 45.376 10.368 ;
  LAYER M1 ;
        RECT 45.408 4.836 45.44 10.368 ;
  LAYER M1 ;
        RECT 45.472 4.836 45.504 10.368 ;
  LAYER M1 ;
        RECT 45.536 4.836 45.568 10.368 ;
  LAYER M1 ;
        RECT 45.6 4.836 45.632 10.368 ;
  LAYER M1 ;
        RECT 45.664 4.836 45.696 10.368 ;
  LAYER M1 ;
        RECT 45.728 4.836 45.76 10.368 ;
  LAYER M1 ;
        RECT 45.792 4.836 45.824 10.368 ;
  LAYER M1 ;
        RECT 45.856 4.836 45.888 10.368 ;
  LAYER M1 ;
        RECT 45.92 4.836 45.952 10.368 ;
  LAYER M1 ;
        RECT 45.984 4.836 46.016 10.368 ;
  LAYER M1 ;
        RECT 46.048 4.836 46.08 10.368 ;
  LAYER M1 ;
        RECT 46.112 4.836 46.144 10.368 ;
  LAYER M1 ;
        RECT 46.176 4.836 46.208 10.368 ;
  LAYER M1 ;
        RECT 46.24 4.836 46.272 10.368 ;
  LAYER M1 ;
        RECT 46.304 4.836 46.336 10.368 ;
  LAYER M1 ;
        RECT 46.368 4.836 46.4 10.368 ;
  LAYER M1 ;
        RECT 46.432 4.836 46.464 10.368 ;
  LAYER M1 ;
        RECT 46.496 4.836 46.528 10.368 ;
  LAYER M1 ;
        RECT 46.56 4.836 46.592 10.368 ;
  LAYER M1 ;
        RECT 46.624 4.836 46.656 10.368 ;
  LAYER M1 ;
        RECT 46.688 4.836 46.72 10.368 ;
  LAYER M1 ;
        RECT 46.752 4.836 46.784 10.368 ;
  LAYER M1 ;
        RECT 46.816 4.836 46.848 10.368 ;
  LAYER M1 ;
        RECT 46.88 4.836 46.912 10.368 ;
  LAYER M1 ;
        RECT 46.944 4.836 46.976 10.368 ;
  LAYER M1 ;
        RECT 47.008 4.836 47.04 10.368 ;
  LAYER M1 ;
        RECT 47.072 4.836 47.104 10.368 ;
  LAYER M1 ;
        RECT 47.136 4.836 47.168 10.368 ;
  LAYER M1 ;
        RECT 47.2 4.836 47.232 10.368 ;
  LAYER M1 ;
        RECT 47.264 4.836 47.296 10.368 ;
  LAYER M1 ;
        RECT 47.328 4.836 47.36 10.368 ;
  LAYER M1 ;
        RECT 47.392 4.836 47.424 10.368 ;
  LAYER M1 ;
        RECT 47.456 4.836 47.488 10.368 ;
  LAYER M1 ;
        RECT 47.52 4.836 47.552 10.368 ;
  LAYER M1 ;
        RECT 47.584 4.836 47.616 10.368 ;
  LAYER M1 ;
        RECT 47.648 4.836 47.68 10.368 ;
  LAYER M1 ;
        RECT 47.712 4.836 47.744 10.368 ;
  LAYER M1 ;
        RECT 47.776 4.836 47.808 10.368 ;
  LAYER M1 ;
        RECT 47.84 4.836 47.872 10.368 ;
  LAYER M1 ;
        RECT 47.904 4.836 47.936 10.368 ;
  LAYER M1 ;
        RECT 47.968 4.836 48 10.368 ;
  LAYER M1 ;
        RECT 48.032 4.836 48.064 10.368 ;
  LAYER M1 ;
        RECT 48.096 4.836 48.128 10.368 ;
  LAYER M1 ;
        RECT 48.16 4.836 48.192 10.368 ;
  LAYER M1 ;
        RECT 48.224 4.836 48.256 10.368 ;
  LAYER M2 ;
        RECT 42.764 4.92 48.276 4.952 ;
  LAYER M2 ;
        RECT 42.764 4.984 48.276 5.016 ;
  LAYER M2 ;
        RECT 42.764 5.048 48.276 5.08 ;
  LAYER M2 ;
        RECT 42.764 5.112 48.276 5.144 ;
  LAYER M2 ;
        RECT 42.764 5.176 48.276 5.208 ;
  LAYER M2 ;
        RECT 42.764 5.24 48.276 5.272 ;
  LAYER M2 ;
        RECT 42.764 5.304 48.276 5.336 ;
  LAYER M2 ;
        RECT 42.764 5.368 48.276 5.4 ;
  LAYER M2 ;
        RECT 42.764 5.432 48.276 5.464 ;
  LAYER M2 ;
        RECT 42.764 5.496 48.276 5.528 ;
  LAYER M2 ;
        RECT 42.764 5.56 48.276 5.592 ;
  LAYER M2 ;
        RECT 42.764 5.624 48.276 5.656 ;
  LAYER M2 ;
        RECT 42.764 5.688 48.276 5.72 ;
  LAYER M2 ;
        RECT 42.764 5.752 48.276 5.784 ;
  LAYER M2 ;
        RECT 42.764 5.816 48.276 5.848 ;
  LAYER M2 ;
        RECT 42.764 5.88 48.276 5.912 ;
  LAYER M2 ;
        RECT 42.764 5.944 48.276 5.976 ;
  LAYER M2 ;
        RECT 42.764 6.008 48.276 6.04 ;
  LAYER M2 ;
        RECT 42.764 6.072 48.276 6.104 ;
  LAYER M2 ;
        RECT 42.764 6.136 48.276 6.168 ;
  LAYER M2 ;
        RECT 42.764 6.2 48.276 6.232 ;
  LAYER M2 ;
        RECT 42.764 6.264 48.276 6.296 ;
  LAYER M2 ;
        RECT 42.764 6.328 48.276 6.36 ;
  LAYER M2 ;
        RECT 42.764 6.392 48.276 6.424 ;
  LAYER M2 ;
        RECT 42.764 6.456 48.276 6.488 ;
  LAYER M2 ;
        RECT 42.764 6.52 48.276 6.552 ;
  LAYER M2 ;
        RECT 42.764 6.584 48.276 6.616 ;
  LAYER M2 ;
        RECT 42.764 6.648 48.276 6.68 ;
  LAYER M2 ;
        RECT 42.764 6.712 48.276 6.744 ;
  LAYER M2 ;
        RECT 42.764 6.776 48.276 6.808 ;
  LAYER M2 ;
        RECT 42.764 6.84 48.276 6.872 ;
  LAYER M2 ;
        RECT 42.764 6.904 48.276 6.936 ;
  LAYER M2 ;
        RECT 42.764 6.968 48.276 7 ;
  LAYER M2 ;
        RECT 42.764 7.032 48.276 7.064 ;
  LAYER M2 ;
        RECT 42.764 7.096 48.276 7.128 ;
  LAYER M2 ;
        RECT 42.764 7.16 48.276 7.192 ;
  LAYER M2 ;
        RECT 42.764 7.224 48.276 7.256 ;
  LAYER M2 ;
        RECT 42.764 7.288 48.276 7.32 ;
  LAYER M2 ;
        RECT 42.764 7.352 48.276 7.384 ;
  LAYER M2 ;
        RECT 42.764 7.416 48.276 7.448 ;
  LAYER M2 ;
        RECT 42.764 7.48 48.276 7.512 ;
  LAYER M2 ;
        RECT 42.764 7.544 48.276 7.576 ;
  LAYER M2 ;
        RECT 42.764 7.608 48.276 7.64 ;
  LAYER M2 ;
        RECT 42.764 7.672 48.276 7.704 ;
  LAYER M2 ;
        RECT 42.764 7.736 48.276 7.768 ;
  LAYER M2 ;
        RECT 42.764 7.8 48.276 7.832 ;
  LAYER M2 ;
        RECT 42.764 7.864 48.276 7.896 ;
  LAYER M2 ;
        RECT 42.764 7.928 48.276 7.96 ;
  LAYER M2 ;
        RECT 42.764 7.992 48.276 8.024 ;
  LAYER M2 ;
        RECT 42.764 8.056 48.276 8.088 ;
  LAYER M2 ;
        RECT 42.764 8.12 48.276 8.152 ;
  LAYER M2 ;
        RECT 42.764 8.184 48.276 8.216 ;
  LAYER M2 ;
        RECT 42.764 8.248 48.276 8.28 ;
  LAYER M2 ;
        RECT 42.764 8.312 48.276 8.344 ;
  LAYER M2 ;
        RECT 42.764 8.376 48.276 8.408 ;
  LAYER M2 ;
        RECT 42.764 8.44 48.276 8.472 ;
  LAYER M2 ;
        RECT 42.764 8.504 48.276 8.536 ;
  LAYER M2 ;
        RECT 42.764 8.568 48.276 8.6 ;
  LAYER M2 ;
        RECT 42.764 8.632 48.276 8.664 ;
  LAYER M2 ;
        RECT 42.764 8.696 48.276 8.728 ;
  LAYER M2 ;
        RECT 42.764 8.76 48.276 8.792 ;
  LAYER M2 ;
        RECT 42.764 8.824 48.276 8.856 ;
  LAYER M2 ;
        RECT 42.764 8.888 48.276 8.92 ;
  LAYER M2 ;
        RECT 42.764 8.952 48.276 8.984 ;
  LAYER M2 ;
        RECT 42.764 9.016 48.276 9.048 ;
  LAYER M2 ;
        RECT 42.764 9.08 48.276 9.112 ;
  LAYER M2 ;
        RECT 42.764 9.144 48.276 9.176 ;
  LAYER M2 ;
        RECT 42.764 9.208 48.276 9.24 ;
  LAYER M2 ;
        RECT 42.764 9.272 48.276 9.304 ;
  LAYER M2 ;
        RECT 42.764 9.336 48.276 9.368 ;
  LAYER M2 ;
        RECT 42.764 9.4 48.276 9.432 ;
  LAYER M2 ;
        RECT 42.764 9.464 48.276 9.496 ;
  LAYER M2 ;
        RECT 42.764 9.528 48.276 9.56 ;
  LAYER M2 ;
        RECT 42.764 9.592 48.276 9.624 ;
  LAYER M2 ;
        RECT 42.764 9.656 48.276 9.688 ;
  LAYER M2 ;
        RECT 42.764 9.72 48.276 9.752 ;
  LAYER M2 ;
        RECT 42.764 9.784 48.276 9.816 ;
  LAYER M2 ;
        RECT 42.764 9.848 48.276 9.88 ;
  LAYER M2 ;
        RECT 42.764 9.912 48.276 9.944 ;
  LAYER M2 ;
        RECT 42.764 9.976 48.276 10.008 ;
  LAYER M2 ;
        RECT 42.764 10.04 48.276 10.072 ;
  LAYER M2 ;
        RECT 42.764 10.104 48.276 10.136 ;
  LAYER M2 ;
        RECT 42.764 10.168 48.276 10.2 ;
  LAYER M2 ;
        RECT 42.764 10.232 48.276 10.264 ;
  LAYER M3 ;
        RECT 42.784 4.836 42.816 10.368 ;
  LAYER M3 ;
        RECT 42.848 4.836 42.88 10.368 ;
  LAYER M3 ;
        RECT 42.912 4.836 42.944 10.368 ;
  LAYER M3 ;
        RECT 42.976 4.836 43.008 10.368 ;
  LAYER M3 ;
        RECT 43.04 4.836 43.072 10.368 ;
  LAYER M3 ;
        RECT 43.104 4.836 43.136 10.368 ;
  LAYER M3 ;
        RECT 43.168 4.836 43.2 10.368 ;
  LAYER M3 ;
        RECT 43.232 4.836 43.264 10.368 ;
  LAYER M3 ;
        RECT 43.296 4.836 43.328 10.368 ;
  LAYER M3 ;
        RECT 43.36 4.836 43.392 10.368 ;
  LAYER M3 ;
        RECT 43.424 4.836 43.456 10.368 ;
  LAYER M3 ;
        RECT 43.488 4.836 43.52 10.368 ;
  LAYER M3 ;
        RECT 43.552 4.836 43.584 10.368 ;
  LAYER M3 ;
        RECT 43.616 4.836 43.648 10.368 ;
  LAYER M3 ;
        RECT 43.68 4.836 43.712 10.368 ;
  LAYER M3 ;
        RECT 43.744 4.836 43.776 10.368 ;
  LAYER M3 ;
        RECT 43.808 4.836 43.84 10.368 ;
  LAYER M3 ;
        RECT 43.872 4.836 43.904 10.368 ;
  LAYER M3 ;
        RECT 43.936 4.836 43.968 10.368 ;
  LAYER M3 ;
        RECT 44 4.836 44.032 10.368 ;
  LAYER M3 ;
        RECT 44.064 4.836 44.096 10.368 ;
  LAYER M3 ;
        RECT 44.128 4.836 44.16 10.368 ;
  LAYER M3 ;
        RECT 44.192 4.836 44.224 10.368 ;
  LAYER M3 ;
        RECT 44.256 4.836 44.288 10.368 ;
  LAYER M3 ;
        RECT 44.32 4.836 44.352 10.368 ;
  LAYER M3 ;
        RECT 44.384 4.836 44.416 10.368 ;
  LAYER M3 ;
        RECT 44.448 4.836 44.48 10.368 ;
  LAYER M3 ;
        RECT 44.512 4.836 44.544 10.368 ;
  LAYER M3 ;
        RECT 44.576 4.836 44.608 10.368 ;
  LAYER M3 ;
        RECT 44.64 4.836 44.672 10.368 ;
  LAYER M3 ;
        RECT 44.704 4.836 44.736 10.368 ;
  LAYER M3 ;
        RECT 44.768 4.836 44.8 10.368 ;
  LAYER M3 ;
        RECT 44.832 4.836 44.864 10.368 ;
  LAYER M3 ;
        RECT 44.896 4.836 44.928 10.368 ;
  LAYER M3 ;
        RECT 44.96 4.836 44.992 10.368 ;
  LAYER M3 ;
        RECT 45.024 4.836 45.056 10.368 ;
  LAYER M3 ;
        RECT 45.088 4.836 45.12 10.368 ;
  LAYER M3 ;
        RECT 45.152 4.836 45.184 10.368 ;
  LAYER M3 ;
        RECT 45.216 4.836 45.248 10.368 ;
  LAYER M3 ;
        RECT 45.28 4.836 45.312 10.368 ;
  LAYER M3 ;
        RECT 45.344 4.836 45.376 10.368 ;
  LAYER M3 ;
        RECT 45.408 4.836 45.44 10.368 ;
  LAYER M3 ;
        RECT 45.472 4.836 45.504 10.368 ;
  LAYER M3 ;
        RECT 45.536 4.836 45.568 10.368 ;
  LAYER M3 ;
        RECT 45.6 4.836 45.632 10.368 ;
  LAYER M3 ;
        RECT 45.664 4.836 45.696 10.368 ;
  LAYER M3 ;
        RECT 45.728 4.836 45.76 10.368 ;
  LAYER M3 ;
        RECT 45.792 4.836 45.824 10.368 ;
  LAYER M3 ;
        RECT 45.856 4.836 45.888 10.368 ;
  LAYER M3 ;
        RECT 45.92 4.836 45.952 10.368 ;
  LAYER M3 ;
        RECT 45.984 4.836 46.016 10.368 ;
  LAYER M3 ;
        RECT 46.048 4.836 46.08 10.368 ;
  LAYER M3 ;
        RECT 46.112 4.836 46.144 10.368 ;
  LAYER M3 ;
        RECT 46.176 4.836 46.208 10.368 ;
  LAYER M3 ;
        RECT 46.24 4.836 46.272 10.368 ;
  LAYER M3 ;
        RECT 46.304 4.836 46.336 10.368 ;
  LAYER M3 ;
        RECT 46.368 4.836 46.4 10.368 ;
  LAYER M3 ;
        RECT 46.432 4.836 46.464 10.368 ;
  LAYER M3 ;
        RECT 46.496 4.836 46.528 10.368 ;
  LAYER M3 ;
        RECT 46.56 4.836 46.592 10.368 ;
  LAYER M3 ;
        RECT 46.624 4.836 46.656 10.368 ;
  LAYER M3 ;
        RECT 46.688 4.836 46.72 10.368 ;
  LAYER M3 ;
        RECT 46.752 4.836 46.784 10.368 ;
  LAYER M3 ;
        RECT 46.816 4.836 46.848 10.368 ;
  LAYER M3 ;
        RECT 46.88 4.836 46.912 10.368 ;
  LAYER M3 ;
        RECT 46.944 4.836 46.976 10.368 ;
  LAYER M3 ;
        RECT 47.008 4.836 47.04 10.368 ;
  LAYER M3 ;
        RECT 47.072 4.836 47.104 10.368 ;
  LAYER M3 ;
        RECT 47.136 4.836 47.168 10.368 ;
  LAYER M3 ;
        RECT 47.2 4.836 47.232 10.368 ;
  LAYER M3 ;
        RECT 47.264 4.836 47.296 10.368 ;
  LAYER M3 ;
        RECT 47.328 4.836 47.36 10.368 ;
  LAYER M3 ;
        RECT 47.392 4.836 47.424 10.368 ;
  LAYER M3 ;
        RECT 47.456 4.836 47.488 10.368 ;
  LAYER M3 ;
        RECT 47.52 4.836 47.552 10.368 ;
  LAYER M3 ;
        RECT 47.584 4.836 47.616 10.368 ;
  LAYER M3 ;
        RECT 47.648 4.836 47.68 10.368 ;
  LAYER M3 ;
        RECT 47.712 4.836 47.744 10.368 ;
  LAYER M3 ;
        RECT 47.776 4.836 47.808 10.368 ;
  LAYER M3 ;
        RECT 47.84 4.836 47.872 10.368 ;
  LAYER M3 ;
        RECT 47.904 4.836 47.936 10.368 ;
  LAYER M3 ;
        RECT 47.968 4.836 48 10.368 ;
  LAYER M3 ;
        RECT 48.032 4.836 48.064 10.368 ;
  LAYER M3 ;
        RECT 48.096 4.836 48.128 10.368 ;
  LAYER M3 ;
        RECT 48.16 4.836 48.192 10.368 ;
  LAYER M3 ;
        RECT 48.22 4.836 48.26 10.368 ;
  LAYER M2 ;
        RECT 42.524 10.316 48.516 10.348 ;
  LAYER M2 ;
        RECT 42.524 4.856 48.516 4.888 ;
  LAYER M1 ;
        RECT 36.704 4.836 36.736 10.368 ;
  LAYER M1 ;
        RECT 36.768 4.836 36.8 10.368 ;
  LAYER M1 ;
        RECT 36.832 4.836 36.864 10.368 ;
  LAYER M1 ;
        RECT 36.896 4.836 36.928 10.368 ;
  LAYER M1 ;
        RECT 36.96 4.836 36.992 10.368 ;
  LAYER M1 ;
        RECT 37.024 4.836 37.056 10.368 ;
  LAYER M1 ;
        RECT 37.088 4.836 37.12 10.368 ;
  LAYER M1 ;
        RECT 37.152 4.836 37.184 10.368 ;
  LAYER M1 ;
        RECT 37.216 4.836 37.248 10.368 ;
  LAYER M1 ;
        RECT 37.28 4.836 37.312 10.368 ;
  LAYER M1 ;
        RECT 37.344 4.836 37.376 10.368 ;
  LAYER M1 ;
        RECT 37.408 4.836 37.44 10.368 ;
  LAYER M1 ;
        RECT 37.472 4.836 37.504 10.368 ;
  LAYER M1 ;
        RECT 37.536 4.836 37.568 10.368 ;
  LAYER M1 ;
        RECT 37.6 4.836 37.632 10.368 ;
  LAYER M1 ;
        RECT 37.664 4.836 37.696 10.368 ;
  LAYER M1 ;
        RECT 37.728 4.836 37.76 10.368 ;
  LAYER M1 ;
        RECT 37.792 4.836 37.824 10.368 ;
  LAYER M1 ;
        RECT 37.856 4.836 37.888 10.368 ;
  LAYER M1 ;
        RECT 37.92 4.836 37.952 10.368 ;
  LAYER M1 ;
        RECT 37.984 4.836 38.016 10.368 ;
  LAYER M1 ;
        RECT 38.048 4.836 38.08 10.368 ;
  LAYER M1 ;
        RECT 38.112 4.836 38.144 10.368 ;
  LAYER M1 ;
        RECT 38.176 4.836 38.208 10.368 ;
  LAYER M1 ;
        RECT 38.24 4.836 38.272 10.368 ;
  LAYER M1 ;
        RECT 38.304 4.836 38.336 10.368 ;
  LAYER M1 ;
        RECT 38.368 4.836 38.4 10.368 ;
  LAYER M1 ;
        RECT 38.432 4.836 38.464 10.368 ;
  LAYER M1 ;
        RECT 38.496 4.836 38.528 10.368 ;
  LAYER M1 ;
        RECT 38.56 4.836 38.592 10.368 ;
  LAYER M1 ;
        RECT 38.624 4.836 38.656 10.368 ;
  LAYER M1 ;
        RECT 38.688 4.836 38.72 10.368 ;
  LAYER M1 ;
        RECT 38.752 4.836 38.784 10.368 ;
  LAYER M1 ;
        RECT 38.816 4.836 38.848 10.368 ;
  LAYER M1 ;
        RECT 38.88 4.836 38.912 10.368 ;
  LAYER M1 ;
        RECT 38.944 4.836 38.976 10.368 ;
  LAYER M1 ;
        RECT 39.008 4.836 39.04 10.368 ;
  LAYER M1 ;
        RECT 39.072 4.836 39.104 10.368 ;
  LAYER M1 ;
        RECT 39.136 4.836 39.168 10.368 ;
  LAYER M1 ;
        RECT 39.2 4.836 39.232 10.368 ;
  LAYER M1 ;
        RECT 39.264 4.836 39.296 10.368 ;
  LAYER M1 ;
        RECT 39.328 4.836 39.36 10.368 ;
  LAYER M1 ;
        RECT 39.392 4.836 39.424 10.368 ;
  LAYER M1 ;
        RECT 39.456 4.836 39.488 10.368 ;
  LAYER M1 ;
        RECT 39.52 4.836 39.552 10.368 ;
  LAYER M1 ;
        RECT 39.584 4.836 39.616 10.368 ;
  LAYER M1 ;
        RECT 39.648 4.836 39.68 10.368 ;
  LAYER M1 ;
        RECT 39.712 4.836 39.744 10.368 ;
  LAYER M1 ;
        RECT 39.776 4.836 39.808 10.368 ;
  LAYER M1 ;
        RECT 39.84 4.836 39.872 10.368 ;
  LAYER M1 ;
        RECT 39.904 4.836 39.936 10.368 ;
  LAYER M1 ;
        RECT 39.968 4.836 40 10.368 ;
  LAYER M1 ;
        RECT 40.032 4.836 40.064 10.368 ;
  LAYER M1 ;
        RECT 40.096 4.836 40.128 10.368 ;
  LAYER M1 ;
        RECT 40.16 4.836 40.192 10.368 ;
  LAYER M1 ;
        RECT 40.224 4.836 40.256 10.368 ;
  LAYER M1 ;
        RECT 40.288 4.836 40.32 10.368 ;
  LAYER M1 ;
        RECT 40.352 4.836 40.384 10.368 ;
  LAYER M1 ;
        RECT 40.416 4.836 40.448 10.368 ;
  LAYER M1 ;
        RECT 40.48 4.836 40.512 10.368 ;
  LAYER M1 ;
        RECT 40.544 4.836 40.576 10.368 ;
  LAYER M1 ;
        RECT 40.608 4.836 40.64 10.368 ;
  LAYER M1 ;
        RECT 40.672 4.836 40.704 10.368 ;
  LAYER M1 ;
        RECT 40.736 4.836 40.768 10.368 ;
  LAYER M1 ;
        RECT 40.8 4.836 40.832 10.368 ;
  LAYER M1 ;
        RECT 40.864 4.836 40.896 10.368 ;
  LAYER M1 ;
        RECT 40.928 4.836 40.96 10.368 ;
  LAYER M1 ;
        RECT 40.992 4.836 41.024 10.368 ;
  LAYER M1 ;
        RECT 41.056 4.836 41.088 10.368 ;
  LAYER M1 ;
        RECT 41.12 4.836 41.152 10.368 ;
  LAYER M1 ;
        RECT 41.184 4.836 41.216 10.368 ;
  LAYER M1 ;
        RECT 41.248 4.836 41.28 10.368 ;
  LAYER M1 ;
        RECT 41.312 4.836 41.344 10.368 ;
  LAYER M1 ;
        RECT 41.376 4.836 41.408 10.368 ;
  LAYER M1 ;
        RECT 41.44 4.836 41.472 10.368 ;
  LAYER M1 ;
        RECT 41.504 4.836 41.536 10.368 ;
  LAYER M1 ;
        RECT 41.568 4.836 41.6 10.368 ;
  LAYER M1 ;
        RECT 41.632 4.836 41.664 10.368 ;
  LAYER M1 ;
        RECT 41.696 4.836 41.728 10.368 ;
  LAYER M1 ;
        RECT 41.76 4.836 41.792 10.368 ;
  LAYER M1 ;
        RECT 41.824 4.836 41.856 10.368 ;
  LAYER M1 ;
        RECT 41.888 4.836 41.92 10.368 ;
  LAYER M1 ;
        RECT 41.952 4.836 41.984 10.368 ;
  LAYER M1 ;
        RECT 42.016 4.836 42.048 10.368 ;
  LAYER M1 ;
        RECT 42.08 4.836 42.112 10.368 ;
  LAYER M1 ;
        RECT 42.144 4.836 42.176 10.368 ;
  LAYER M2 ;
        RECT 36.684 4.92 42.196 4.952 ;
  LAYER M2 ;
        RECT 36.684 4.984 42.196 5.016 ;
  LAYER M2 ;
        RECT 36.684 5.048 42.196 5.08 ;
  LAYER M2 ;
        RECT 36.684 5.112 42.196 5.144 ;
  LAYER M2 ;
        RECT 36.684 5.176 42.196 5.208 ;
  LAYER M2 ;
        RECT 36.684 5.24 42.196 5.272 ;
  LAYER M2 ;
        RECT 36.684 5.304 42.196 5.336 ;
  LAYER M2 ;
        RECT 36.684 5.368 42.196 5.4 ;
  LAYER M2 ;
        RECT 36.684 5.432 42.196 5.464 ;
  LAYER M2 ;
        RECT 36.684 5.496 42.196 5.528 ;
  LAYER M2 ;
        RECT 36.684 5.56 42.196 5.592 ;
  LAYER M2 ;
        RECT 36.684 5.624 42.196 5.656 ;
  LAYER M2 ;
        RECT 36.684 5.688 42.196 5.72 ;
  LAYER M2 ;
        RECT 36.684 5.752 42.196 5.784 ;
  LAYER M2 ;
        RECT 36.684 5.816 42.196 5.848 ;
  LAYER M2 ;
        RECT 36.684 5.88 42.196 5.912 ;
  LAYER M2 ;
        RECT 36.684 5.944 42.196 5.976 ;
  LAYER M2 ;
        RECT 36.684 6.008 42.196 6.04 ;
  LAYER M2 ;
        RECT 36.684 6.072 42.196 6.104 ;
  LAYER M2 ;
        RECT 36.684 6.136 42.196 6.168 ;
  LAYER M2 ;
        RECT 36.684 6.2 42.196 6.232 ;
  LAYER M2 ;
        RECT 36.684 6.264 42.196 6.296 ;
  LAYER M2 ;
        RECT 36.684 6.328 42.196 6.36 ;
  LAYER M2 ;
        RECT 36.684 6.392 42.196 6.424 ;
  LAYER M2 ;
        RECT 36.684 6.456 42.196 6.488 ;
  LAYER M2 ;
        RECT 36.684 6.52 42.196 6.552 ;
  LAYER M2 ;
        RECT 36.684 6.584 42.196 6.616 ;
  LAYER M2 ;
        RECT 36.684 6.648 42.196 6.68 ;
  LAYER M2 ;
        RECT 36.684 6.712 42.196 6.744 ;
  LAYER M2 ;
        RECT 36.684 6.776 42.196 6.808 ;
  LAYER M2 ;
        RECT 36.684 6.84 42.196 6.872 ;
  LAYER M2 ;
        RECT 36.684 6.904 42.196 6.936 ;
  LAYER M2 ;
        RECT 36.684 6.968 42.196 7 ;
  LAYER M2 ;
        RECT 36.684 7.032 42.196 7.064 ;
  LAYER M2 ;
        RECT 36.684 7.096 42.196 7.128 ;
  LAYER M2 ;
        RECT 36.684 7.16 42.196 7.192 ;
  LAYER M2 ;
        RECT 36.684 7.224 42.196 7.256 ;
  LAYER M2 ;
        RECT 36.684 7.288 42.196 7.32 ;
  LAYER M2 ;
        RECT 36.684 7.352 42.196 7.384 ;
  LAYER M2 ;
        RECT 36.684 7.416 42.196 7.448 ;
  LAYER M2 ;
        RECT 36.684 7.48 42.196 7.512 ;
  LAYER M2 ;
        RECT 36.684 7.544 42.196 7.576 ;
  LAYER M2 ;
        RECT 36.684 7.608 42.196 7.64 ;
  LAYER M2 ;
        RECT 36.684 7.672 42.196 7.704 ;
  LAYER M2 ;
        RECT 36.684 7.736 42.196 7.768 ;
  LAYER M2 ;
        RECT 36.684 7.8 42.196 7.832 ;
  LAYER M2 ;
        RECT 36.684 7.864 42.196 7.896 ;
  LAYER M2 ;
        RECT 36.684 7.928 42.196 7.96 ;
  LAYER M2 ;
        RECT 36.684 7.992 42.196 8.024 ;
  LAYER M2 ;
        RECT 36.684 8.056 42.196 8.088 ;
  LAYER M2 ;
        RECT 36.684 8.12 42.196 8.152 ;
  LAYER M2 ;
        RECT 36.684 8.184 42.196 8.216 ;
  LAYER M2 ;
        RECT 36.684 8.248 42.196 8.28 ;
  LAYER M2 ;
        RECT 36.684 8.312 42.196 8.344 ;
  LAYER M2 ;
        RECT 36.684 8.376 42.196 8.408 ;
  LAYER M2 ;
        RECT 36.684 8.44 42.196 8.472 ;
  LAYER M2 ;
        RECT 36.684 8.504 42.196 8.536 ;
  LAYER M2 ;
        RECT 36.684 8.568 42.196 8.6 ;
  LAYER M2 ;
        RECT 36.684 8.632 42.196 8.664 ;
  LAYER M2 ;
        RECT 36.684 8.696 42.196 8.728 ;
  LAYER M2 ;
        RECT 36.684 8.76 42.196 8.792 ;
  LAYER M2 ;
        RECT 36.684 8.824 42.196 8.856 ;
  LAYER M2 ;
        RECT 36.684 8.888 42.196 8.92 ;
  LAYER M2 ;
        RECT 36.684 8.952 42.196 8.984 ;
  LAYER M2 ;
        RECT 36.684 9.016 42.196 9.048 ;
  LAYER M2 ;
        RECT 36.684 9.08 42.196 9.112 ;
  LAYER M2 ;
        RECT 36.684 9.144 42.196 9.176 ;
  LAYER M2 ;
        RECT 36.684 9.208 42.196 9.24 ;
  LAYER M2 ;
        RECT 36.684 9.272 42.196 9.304 ;
  LAYER M2 ;
        RECT 36.684 9.336 42.196 9.368 ;
  LAYER M2 ;
        RECT 36.684 9.4 42.196 9.432 ;
  LAYER M2 ;
        RECT 36.684 9.464 42.196 9.496 ;
  LAYER M2 ;
        RECT 36.684 9.528 42.196 9.56 ;
  LAYER M2 ;
        RECT 36.684 9.592 42.196 9.624 ;
  LAYER M2 ;
        RECT 36.684 9.656 42.196 9.688 ;
  LAYER M2 ;
        RECT 36.684 9.72 42.196 9.752 ;
  LAYER M2 ;
        RECT 36.684 9.784 42.196 9.816 ;
  LAYER M2 ;
        RECT 36.684 9.848 42.196 9.88 ;
  LAYER M2 ;
        RECT 36.684 9.912 42.196 9.944 ;
  LAYER M2 ;
        RECT 36.684 9.976 42.196 10.008 ;
  LAYER M2 ;
        RECT 36.684 10.04 42.196 10.072 ;
  LAYER M2 ;
        RECT 36.684 10.104 42.196 10.136 ;
  LAYER M2 ;
        RECT 36.684 10.168 42.196 10.2 ;
  LAYER M2 ;
        RECT 36.684 10.232 42.196 10.264 ;
  LAYER M3 ;
        RECT 36.704 4.836 36.736 10.368 ;
  LAYER M3 ;
        RECT 36.768 4.836 36.8 10.368 ;
  LAYER M3 ;
        RECT 36.832 4.836 36.864 10.368 ;
  LAYER M3 ;
        RECT 36.896 4.836 36.928 10.368 ;
  LAYER M3 ;
        RECT 36.96 4.836 36.992 10.368 ;
  LAYER M3 ;
        RECT 37.024 4.836 37.056 10.368 ;
  LAYER M3 ;
        RECT 37.088 4.836 37.12 10.368 ;
  LAYER M3 ;
        RECT 37.152 4.836 37.184 10.368 ;
  LAYER M3 ;
        RECT 37.216 4.836 37.248 10.368 ;
  LAYER M3 ;
        RECT 37.28 4.836 37.312 10.368 ;
  LAYER M3 ;
        RECT 37.344 4.836 37.376 10.368 ;
  LAYER M3 ;
        RECT 37.408 4.836 37.44 10.368 ;
  LAYER M3 ;
        RECT 37.472 4.836 37.504 10.368 ;
  LAYER M3 ;
        RECT 37.536 4.836 37.568 10.368 ;
  LAYER M3 ;
        RECT 37.6 4.836 37.632 10.368 ;
  LAYER M3 ;
        RECT 37.664 4.836 37.696 10.368 ;
  LAYER M3 ;
        RECT 37.728 4.836 37.76 10.368 ;
  LAYER M3 ;
        RECT 37.792 4.836 37.824 10.368 ;
  LAYER M3 ;
        RECT 37.856 4.836 37.888 10.368 ;
  LAYER M3 ;
        RECT 37.92 4.836 37.952 10.368 ;
  LAYER M3 ;
        RECT 37.984 4.836 38.016 10.368 ;
  LAYER M3 ;
        RECT 38.048 4.836 38.08 10.368 ;
  LAYER M3 ;
        RECT 38.112 4.836 38.144 10.368 ;
  LAYER M3 ;
        RECT 38.176 4.836 38.208 10.368 ;
  LAYER M3 ;
        RECT 38.24 4.836 38.272 10.368 ;
  LAYER M3 ;
        RECT 38.304 4.836 38.336 10.368 ;
  LAYER M3 ;
        RECT 38.368 4.836 38.4 10.368 ;
  LAYER M3 ;
        RECT 38.432 4.836 38.464 10.368 ;
  LAYER M3 ;
        RECT 38.496 4.836 38.528 10.368 ;
  LAYER M3 ;
        RECT 38.56 4.836 38.592 10.368 ;
  LAYER M3 ;
        RECT 38.624 4.836 38.656 10.368 ;
  LAYER M3 ;
        RECT 38.688 4.836 38.72 10.368 ;
  LAYER M3 ;
        RECT 38.752 4.836 38.784 10.368 ;
  LAYER M3 ;
        RECT 38.816 4.836 38.848 10.368 ;
  LAYER M3 ;
        RECT 38.88 4.836 38.912 10.368 ;
  LAYER M3 ;
        RECT 38.944 4.836 38.976 10.368 ;
  LAYER M3 ;
        RECT 39.008 4.836 39.04 10.368 ;
  LAYER M3 ;
        RECT 39.072 4.836 39.104 10.368 ;
  LAYER M3 ;
        RECT 39.136 4.836 39.168 10.368 ;
  LAYER M3 ;
        RECT 39.2 4.836 39.232 10.368 ;
  LAYER M3 ;
        RECT 39.264 4.836 39.296 10.368 ;
  LAYER M3 ;
        RECT 39.328 4.836 39.36 10.368 ;
  LAYER M3 ;
        RECT 39.392 4.836 39.424 10.368 ;
  LAYER M3 ;
        RECT 39.456 4.836 39.488 10.368 ;
  LAYER M3 ;
        RECT 39.52 4.836 39.552 10.368 ;
  LAYER M3 ;
        RECT 39.584 4.836 39.616 10.368 ;
  LAYER M3 ;
        RECT 39.648 4.836 39.68 10.368 ;
  LAYER M3 ;
        RECT 39.712 4.836 39.744 10.368 ;
  LAYER M3 ;
        RECT 39.776 4.836 39.808 10.368 ;
  LAYER M3 ;
        RECT 39.84 4.836 39.872 10.368 ;
  LAYER M3 ;
        RECT 39.904 4.836 39.936 10.368 ;
  LAYER M3 ;
        RECT 39.968 4.836 40 10.368 ;
  LAYER M3 ;
        RECT 40.032 4.836 40.064 10.368 ;
  LAYER M3 ;
        RECT 40.096 4.836 40.128 10.368 ;
  LAYER M3 ;
        RECT 40.16 4.836 40.192 10.368 ;
  LAYER M3 ;
        RECT 40.224 4.836 40.256 10.368 ;
  LAYER M3 ;
        RECT 40.288 4.836 40.32 10.368 ;
  LAYER M3 ;
        RECT 40.352 4.836 40.384 10.368 ;
  LAYER M3 ;
        RECT 40.416 4.836 40.448 10.368 ;
  LAYER M3 ;
        RECT 40.48 4.836 40.512 10.368 ;
  LAYER M3 ;
        RECT 40.544 4.836 40.576 10.368 ;
  LAYER M3 ;
        RECT 40.608 4.836 40.64 10.368 ;
  LAYER M3 ;
        RECT 40.672 4.836 40.704 10.368 ;
  LAYER M3 ;
        RECT 40.736 4.836 40.768 10.368 ;
  LAYER M3 ;
        RECT 40.8 4.836 40.832 10.368 ;
  LAYER M3 ;
        RECT 40.864 4.836 40.896 10.368 ;
  LAYER M3 ;
        RECT 40.928 4.836 40.96 10.368 ;
  LAYER M3 ;
        RECT 40.992 4.836 41.024 10.368 ;
  LAYER M3 ;
        RECT 41.056 4.836 41.088 10.368 ;
  LAYER M3 ;
        RECT 41.12 4.836 41.152 10.368 ;
  LAYER M3 ;
        RECT 41.184 4.836 41.216 10.368 ;
  LAYER M3 ;
        RECT 41.248 4.836 41.28 10.368 ;
  LAYER M3 ;
        RECT 41.312 4.836 41.344 10.368 ;
  LAYER M3 ;
        RECT 41.376 4.836 41.408 10.368 ;
  LAYER M3 ;
        RECT 41.44 4.836 41.472 10.368 ;
  LAYER M3 ;
        RECT 41.504 4.836 41.536 10.368 ;
  LAYER M3 ;
        RECT 41.568 4.836 41.6 10.368 ;
  LAYER M3 ;
        RECT 41.632 4.836 41.664 10.368 ;
  LAYER M3 ;
        RECT 41.696 4.836 41.728 10.368 ;
  LAYER M3 ;
        RECT 41.76 4.836 41.792 10.368 ;
  LAYER M3 ;
        RECT 41.824 4.836 41.856 10.368 ;
  LAYER M3 ;
        RECT 41.888 4.836 41.92 10.368 ;
  LAYER M3 ;
        RECT 41.952 4.836 41.984 10.368 ;
  LAYER M3 ;
        RECT 42.016 4.836 42.048 10.368 ;
  LAYER M3 ;
        RECT 42.08 4.836 42.112 10.368 ;
  LAYER M3 ;
        RECT 42.14 4.836 42.18 10.368 ;
  LAYER M2 ;
        RECT 36.444 10.316 42.436 10.348 ;
  LAYER M2 ;
        RECT 36.444 4.856 42.436 4.888 ;
  LAYER M1 ;
        RECT 15.744 4.836 15.776 10.368 ;
  LAYER M1 ;
        RECT 15.68 4.836 15.712 10.368 ;
  LAYER M1 ;
        RECT 15.616 4.836 15.648 10.368 ;
  LAYER M1 ;
        RECT 15.552 4.836 15.584 10.368 ;
  LAYER M1 ;
        RECT 15.488 4.836 15.52 10.368 ;
  LAYER M1 ;
        RECT 15.424 4.836 15.456 10.368 ;
  LAYER M1 ;
        RECT 15.36 4.836 15.392 10.368 ;
  LAYER M1 ;
        RECT 15.296 4.836 15.328 10.368 ;
  LAYER M1 ;
        RECT 15.232 4.836 15.264 10.368 ;
  LAYER M1 ;
        RECT 15.168 4.836 15.2 10.368 ;
  LAYER M1 ;
        RECT 15.104 4.836 15.136 10.368 ;
  LAYER M1 ;
        RECT 15.04 4.836 15.072 10.368 ;
  LAYER M1 ;
        RECT 14.976 4.836 15.008 10.368 ;
  LAYER M1 ;
        RECT 14.912 4.836 14.944 10.368 ;
  LAYER M1 ;
        RECT 14.848 4.836 14.88 10.368 ;
  LAYER M1 ;
        RECT 14.784 4.836 14.816 10.368 ;
  LAYER M1 ;
        RECT 14.72 4.836 14.752 10.368 ;
  LAYER M1 ;
        RECT 14.656 4.836 14.688 10.368 ;
  LAYER M1 ;
        RECT 14.592 4.836 14.624 10.368 ;
  LAYER M1 ;
        RECT 14.528 4.836 14.56 10.368 ;
  LAYER M1 ;
        RECT 14.464 4.836 14.496 10.368 ;
  LAYER M1 ;
        RECT 14.4 4.836 14.432 10.368 ;
  LAYER M1 ;
        RECT 14.336 4.836 14.368 10.368 ;
  LAYER M1 ;
        RECT 14.272 4.836 14.304 10.368 ;
  LAYER M1 ;
        RECT 14.208 4.836 14.24 10.368 ;
  LAYER M1 ;
        RECT 14.144 4.836 14.176 10.368 ;
  LAYER M1 ;
        RECT 14.08 4.836 14.112 10.368 ;
  LAYER M1 ;
        RECT 14.016 4.836 14.048 10.368 ;
  LAYER M1 ;
        RECT 13.952 4.836 13.984 10.368 ;
  LAYER M1 ;
        RECT 13.888 4.836 13.92 10.368 ;
  LAYER M1 ;
        RECT 13.824 4.836 13.856 10.368 ;
  LAYER M1 ;
        RECT 13.76 4.836 13.792 10.368 ;
  LAYER M1 ;
        RECT 13.696 4.836 13.728 10.368 ;
  LAYER M1 ;
        RECT 13.632 4.836 13.664 10.368 ;
  LAYER M1 ;
        RECT 13.568 4.836 13.6 10.368 ;
  LAYER M1 ;
        RECT 13.504 4.836 13.536 10.368 ;
  LAYER M1 ;
        RECT 13.44 4.836 13.472 10.368 ;
  LAYER M1 ;
        RECT 13.376 4.836 13.408 10.368 ;
  LAYER M1 ;
        RECT 13.312 4.836 13.344 10.368 ;
  LAYER M1 ;
        RECT 13.248 4.836 13.28 10.368 ;
  LAYER M1 ;
        RECT 13.184 4.836 13.216 10.368 ;
  LAYER M1 ;
        RECT 13.12 4.836 13.152 10.368 ;
  LAYER M1 ;
        RECT 13.056 4.836 13.088 10.368 ;
  LAYER M1 ;
        RECT 12.992 4.836 13.024 10.368 ;
  LAYER M1 ;
        RECT 12.928 4.836 12.96 10.368 ;
  LAYER M1 ;
        RECT 12.864 4.836 12.896 10.368 ;
  LAYER M1 ;
        RECT 12.8 4.836 12.832 10.368 ;
  LAYER M1 ;
        RECT 12.736 4.836 12.768 10.368 ;
  LAYER M1 ;
        RECT 12.672 4.836 12.704 10.368 ;
  LAYER M1 ;
        RECT 12.608 4.836 12.64 10.368 ;
  LAYER M1 ;
        RECT 12.544 4.836 12.576 10.368 ;
  LAYER M1 ;
        RECT 12.48 4.836 12.512 10.368 ;
  LAYER M1 ;
        RECT 12.416 4.836 12.448 10.368 ;
  LAYER M1 ;
        RECT 12.352 4.836 12.384 10.368 ;
  LAYER M1 ;
        RECT 12.288 4.836 12.32 10.368 ;
  LAYER M1 ;
        RECT 12.224 4.836 12.256 10.368 ;
  LAYER M1 ;
        RECT 12.16 4.836 12.192 10.368 ;
  LAYER M1 ;
        RECT 12.096 4.836 12.128 10.368 ;
  LAYER M1 ;
        RECT 12.032 4.836 12.064 10.368 ;
  LAYER M1 ;
        RECT 11.968 4.836 12 10.368 ;
  LAYER M1 ;
        RECT 11.904 4.836 11.936 10.368 ;
  LAYER M1 ;
        RECT 11.84 4.836 11.872 10.368 ;
  LAYER M1 ;
        RECT 11.776 4.836 11.808 10.368 ;
  LAYER M1 ;
        RECT 11.712 4.836 11.744 10.368 ;
  LAYER M1 ;
        RECT 11.648 4.836 11.68 10.368 ;
  LAYER M1 ;
        RECT 11.584 4.836 11.616 10.368 ;
  LAYER M1 ;
        RECT 11.52 4.836 11.552 10.368 ;
  LAYER M1 ;
        RECT 11.456 4.836 11.488 10.368 ;
  LAYER M1 ;
        RECT 11.392 4.836 11.424 10.368 ;
  LAYER M1 ;
        RECT 11.328 4.836 11.36 10.368 ;
  LAYER M1 ;
        RECT 11.264 4.836 11.296 10.368 ;
  LAYER M1 ;
        RECT 11.2 4.836 11.232 10.368 ;
  LAYER M1 ;
        RECT 11.136 4.836 11.168 10.368 ;
  LAYER M1 ;
        RECT 11.072 4.836 11.104 10.368 ;
  LAYER M1 ;
        RECT 11.008 4.836 11.04 10.368 ;
  LAYER M1 ;
        RECT 10.944 4.836 10.976 10.368 ;
  LAYER M1 ;
        RECT 10.88 4.836 10.912 10.368 ;
  LAYER M1 ;
        RECT 10.816 4.836 10.848 10.368 ;
  LAYER M1 ;
        RECT 10.752 4.836 10.784 10.368 ;
  LAYER M1 ;
        RECT 10.688 4.836 10.72 10.368 ;
  LAYER M1 ;
        RECT 10.624 4.836 10.656 10.368 ;
  LAYER M1 ;
        RECT 10.56 4.836 10.592 10.368 ;
  LAYER M1 ;
        RECT 10.496 4.836 10.528 10.368 ;
  LAYER M1 ;
        RECT 10.432 4.836 10.464 10.368 ;
  LAYER M1 ;
        RECT 10.368 4.836 10.4 10.368 ;
  LAYER M1 ;
        RECT 10.304 4.836 10.336 10.368 ;
  LAYER M2 ;
        RECT 10.284 4.92 15.796 4.952 ;
  LAYER M2 ;
        RECT 10.284 4.984 15.796 5.016 ;
  LAYER M2 ;
        RECT 10.284 5.048 15.796 5.08 ;
  LAYER M2 ;
        RECT 10.284 5.112 15.796 5.144 ;
  LAYER M2 ;
        RECT 10.284 5.176 15.796 5.208 ;
  LAYER M2 ;
        RECT 10.284 5.24 15.796 5.272 ;
  LAYER M2 ;
        RECT 10.284 5.304 15.796 5.336 ;
  LAYER M2 ;
        RECT 10.284 5.368 15.796 5.4 ;
  LAYER M2 ;
        RECT 10.284 5.432 15.796 5.464 ;
  LAYER M2 ;
        RECT 10.284 5.496 15.796 5.528 ;
  LAYER M2 ;
        RECT 10.284 5.56 15.796 5.592 ;
  LAYER M2 ;
        RECT 10.284 5.624 15.796 5.656 ;
  LAYER M2 ;
        RECT 10.284 5.688 15.796 5.72 ;
  LAYER M2 ;
        RECT 10.284 5.752 15.796 5.784 ;
  LAYER M2 ;
        RECT 10.284 5.816 15.796 5.848 ;
  LAYER M2 ;
        RECT 10.284 5.88 15.796 5.912 ;
  LAYER M2 ;
        RECT 10.284 5.944 15.796 5.976 ;
  LAYER M2 ;
        RECT 10.284 6.008 15.796 6.04 ;
  LAYER M2 ;
        RECT 10.284 6.072 15.796 6.104 ;
  LAYER M2 ;
        RECT 10.284 6.136 15.796 6.168 ;
  LAYER M2 ;
        RECT 10.284 6.2 15.796 6.232 ;
  LAYER M2 ;
        RECT 10.284 6.264 15.796 6.296 ;
  LAYER M2 ;
        RECT 10.284 6.328 15.796 6.36 ;
  LAYER M2 ;
        RECT 10.284 6.392 15.796 6.424 ;
  LAYER M2 ;
        RECT 10.284 6.456 15.796 6.488 ;
  LAYER M2 ;
        RECT 10.284 6.52 15.796 6.552 ;
  LAYER M2 ;
        RECT 10.284 6.584 15.796 6.616 ;
  LAYER M2 ;
        RECT 10.284 6.648 15.796 6.68 ;
  LAYER M2 ;
        RECT 10.284 6.712 15.796 6.744 ;
  LAYER M2 ;
        RECT 10.284 6.776 15.796 6.808 ;
  LAYER M2 ;
        RECT 10.284 6.84 15.796 6.872 ;
  LAYER M2 ;
        RECT 10.284 6.904 15.796 6.936 ;
  LAYER M2 ;
        RECT 10.284 6.968 15.796 7 ;
  LAYER M2 ;
        RECT 10.284 7.032 15.796 7.064 ;
  LAYER M2 ;
        RECT 10.284 7.096 15.796 7.128 ;
  LAYER M2 ;
        RECT 10.284 7.16 15.796 7.192 ;
  LAYER M2 ;
        RECT 10.284 7.224 15.796 7.256 ;
  LAYER M2 ;
        RECT 10.284 7.288 15.796 7.32 ;
  LAYER M2 ;
        RECT 10.284 7.352 15.796 7.384 ;
  LAYER M2 ;
        RECT 10.284 7.416 15.796 7.448 ;
  LAYER M2 ;
        RECT 10.284 7.48 15.796 7.512 ;
  LAYER M2 ;
        RECT 10.284 7.544 15.796 7.576 ;
  LAYER M2 ;
        RECT 10.284 7.608 15.796 7.64 ;
  LAYER M2 ;
        RECT 10.284 7.672 15.796 7.704 ;
  LAYER M2 ;
        RECT 10.284 7.736 15.796 7.768 ;
  LAYER M2 ;
        RECT 10.284 7.8 15.796 7.832 ;
  LAYER M2 ;
        RECT 10.284 7.864 15.796 7.896 ;
  LAYER M2 ;
        RECT 10.284 7.928 15.796 7.96 ;
  LAYER M2 ;
        RECT 10.284 7.992 15.796 8.024 ;
  LAYER M2 ;
        RECT 10.284 8.056 15.796 8.088 ;
  LAYER M2 ;
        RECT 10.284 8.12 15.796 8.152 ;
  LAYER M2 ;
        RECT 10.284 8.184 15.796 8.216 ;
  LAYER M2 ;
        RECT 10.284 8.248 15.796 8.28 ;
  LAYER M2 ;
        RECT 10.284 8.312 15.796 8.344 ;
  LAYER M2 ;
        RECT 10.284 8.376 15.796 8.408 ;
  LAYER M2 ;
        RECT 10.284 8.44 15.796 8.472 ;
  LAYER M2 ;
        RECT 10.284 8.504 15.796 8.536 ;
  LAYER M2 ;
        RECT 10.284 8.568 15.796 8.6 ;
  LAYER M2 ;
        RECT 10.284 8.632 15.796 8.664 ;
  LAYER M2 ;
        RECT 10.284 8.696 15.796 8.728 ;
  LAYER M2 ;
        RECT 10.284 8.76 15.796 8.792 ;
  LAYER M2 ;
        RECT 10.284 8.824 15.796 8.856 ;
  LAYER M2 ;
        RECT 10.284 8.888 15.796 8.92 ;
  LAYER M2 ;
        RECT 10.284 8.952 15.796 8.984 ;
  LAYER M2 ;
        RECT 10.284 9.016 15.796 9.048 ;
  LAYER M2 ;
        RECT 10.284 9.08 15.796 9.112 ;
  LAYER M2 ;
        RECT 10.284 9.144 15.796 9.176 ;
  LAYER M2 ;
        RECT 10.284 9.208 15.796 9.24 ;
  LAYER M2 ;
        RECT 10.284 9.272 15.796 9.304 ;
  LAYER M2 ;
        RECT 10.284 9.336 15.796 9.368 ;
  LAYER M2 ;
        RECT 10.284 9.4 15.796 9.432 ;
  LAYER M2 ;
        RECT 10.284 9.464 15.796 9.496 ;
  LAYER M2 ;
        RECT 10.284 9.528 15.796 9.56 ;
  LAYER M2 ;
        RECT 10.284 9.592 15.796 9.624 ;
  LAYER M2 ;
        RECT 10.284 9.656 15.796 9.688 ;
  LAYER M2 ;
        RECT 10.284 9.72 15.796 9.752 ;
  LAYER M2 ;
        RECT 10.284 9.784 15.796 9.816 ;
  LAYER M2 ;
        RECT 10.284 9.848 15.796 9.88 ;
  LAYER M2 ;
        RECT 10.284 9.912 15.796 9.944 ;
  LAYER M2 ;
        RECT 10.284 9.976 15.796 10.008 ;
  LAYER M2 ;
        RECT 10.284 10.04 15.796 10.072 ;
  LAYER M2 ;
        RECT 10.284 10.104 15.796 10.136 ;
  LAYER M2 ;
        RECT 10.284 10.168 15.796 10.2 ;
  LAYER M2 ;
        RECT 10.284 10.232 15.796 10.264 ;
  LAYER M3 ;
        RECT 15.744 4.836 15.776 10.368 ;
  LAYER M3 ;
        RECT 15.68 4.836 15.712 10.368 ;
  LAYER M3 ;
        RECT 15.616 4.836 15.648 10.368 ;
  LAYER M3 ;
        RECT 15.552 4.836 15.584 10.368 ;
  LAYER M3 ;
        RECT 15.488 4.836 15.52 10.368 ;
  LAYER M3 ;
        RECT 15.424 4.836 15.456 10.368 ;
  LAYER M3 ;
        RECT 15.36 4.836 15.392 10.368 ;
  LAYER M3 ;
        RECT 15.296 4.836 15.328 10.368 ;
  LAYER M3 ;
        RECT 15.232 4.836 15.264 10.368 ;
  LAYER M3 ;
        RECT 15.168 4.836 15.2 10.368 ;
  LAYER M3 ;
        RECT 15.104 4.836 15.136 10.368 ;
  LAYER M3 ;
        RECT 15.04 4.836 15.072 10.368 ;
  LAYER M3 ;
        RECT 14.976 4.836 15.008 10.368 ;
  LAYER M3 ;
        RECT 14.912 4.836 14.944 10.368 ;
  LAYER M3 ;
        RECT 14.848 4.836 14.88 10.368 ;
  LAYER M3 ;
        RECT 14.784 4.836 14.816 10.368 ;
  LAYER M3 ;
        RECT 14.72 4.836 14.752 10.368 ;
  LAYER M3 ;
        RECT 14.656 4.836 14.688 10.368 ;
  LAYER M3 ;
        RECT 14.592 4.836 14.624 10.368 ;
  LAYER M3 ;
        RECT 14.528 4.836 14.56 10.368 ;
  LAYER M3 ;
        RECT 14.464 4.836 14.496 10.368 ;
  LAYER M3 ;
        RECT 14.4 4.836 14.432 10.368 ;
  LAYER M3 ;
        RECT 14.336 4.836 14.368 10.368 ;
  LAYER M3 ;
        RECT 14.272 4.836 14.304 10.368 ;
  LAYER M3 ;
        RECT 14.208 4.836 14.24 10.368 ;
  LAYER M3 ;
        RECT 14.144 4.836 14.176 10.368 ;
  LAYER M3 ;
        RECT 14.08 4.836 14.112 10.368 ;
  LAYER M3 ;
        RECT 14.016 4.836 14.048 10.368 ;
  LAYER M3 ;
        RECT 13.952 4.836 13.984 10.368 ;
  LAYER M3 ;
        RECT 13.888 4.836 13.92 10.368 ;
  LAYER M3 ;
        RECT 13.824 4.836 13.856 10.368 ;
  LAYER M3 ;
        RECT 13.76 4.836 13.792 10.368 ;
  LAYER M3 ;
        RECT 13.696 4.836 13.728 10.368 ;
  LAYER M3 ;
        RECT 13.632 4.836 13.664 10.368 ;
  LAYER M3 ;
        RECT 13.568 4.836 13.6 10.368 ;
  LAYER M3 ;
        RECT 13.504 4.836 13.536 10.368 ;
  LAYER M3 ;
        RECT 13.44 4.836 13.472 10.368 ;
  LAYER M3 ;
        RECT 13.376 4.836 13.408 10.368 ;
  LAYER M3 ;
        RECT 13.312 4.836 13.344 10.368 ;
  LAYER M3 ;
        RECT 13.248 4.836 13.28 10.368 ;
  LAYER M3 ;
        RECT 13.184 4.836 13.216 10.368 ;
  LAYER M3 ;
        RECT 13.12 4.836 13.152 10.368 ;
  LAYER M3 ;
        RECT 13.056 4.836 13.088 10.368 ;
  LAYER M3 ;
        RECT 12.992 4.836 13.024 10.368 ;
  LAYER M3 ;
        RECT 12.928 4.836 12.96 10.368 ;
  LAYER M3 ;
        RECT 12.864 4.836 12.896 10.368 ;
  LAYER M3 ;
        RECT 12.8 4.836 12.832 10.368 ;
  LAYER M3 ;
        RECT 12.736 4.836 12.768 10.368 ;
  LAYER M3 ;
        RECT 12.672 4.836 12.704 10.368 ;
  LAYER M3 ;
        RECT 12.608 4.836 12.64 10.368 ;
  LAYER M3 ;
        RECT 12.544 4.836 12.576 10.368 ;
  LAYER M3 ;
        RECT 12.48 4.836 12.512 10.368 ;
  LAYER M3 ;
        RECT 12.416 4.836 12.448 10.368 ;
  LAYER M3 ;
        RECT 12.352 4.836 12.384 10.368 ;
  LAYER M3 ;
        RECT 12.288 4.836 12.32 10.368 ;
  LAYER M3 ;
        RECT 12.224 4.836 12.256 10.368 ;
  LAYER M3 ;
        RECT 12.16 4.836 12.192 10.368 ;
  LAYER M3 ;
        RECT 12.096 4.836 12.128 10.368 ;
  LAYER M3 ;
        RECT 12.032 4.836 12.064 10.368 ;
  LAYER M3 ;
        RECT 11.968 4.836 12 10.368 ;
  LAYER M3 ;
        RECT 11.904 4.836 11.936 10.368 ;
  LAYER M3 ;
        RECT 11.84 4.836 11.872 10.368 ;
  LAYER M3 ;
        RECT 11.776 4.836 11.808 10.368 ;
  LAYER M3 ;
        RECT 11.712 4.836 11.744 10.368 ;
  LAYER M3 ;
        RECT 11.648 4.836 11.68 10.368 ;
  LAYER M3 ;
        RECT 11.584 4.836 11.616 10.368 ;
  LAYER M3 ;
        RECT 11.52 4.836 11.552 10.368 ;
  LAYER M3 ;
        RECT 11.456 4.836 11.488 10.368 ;
  LAYER M3 ;
        RECT 11.392 4.836 11.424 10.368 ;
  LAYER M3 ;
        RECT 11.328 4.836 11.36 10.368 ;
  LAYER M3 ;
        RECT 11.264 4.836 11.296 10.368 ;
  LAYER M3 ;
        RECT 11.2 4.836 11.232 10.368 ;
  LAYER M3 ;
        RECT 11.136 4.836 11.168 10.368 ;
  LAYER M3 ;
        RECT 11.072 4.836 11.104 10.368 ;
  LAYER M3 ;
        RECT 11.008 4.836 11.04 10.368 ;
  LAYER M3 ;
        RECT 10.944 4.836 10.976 10.368 ;
  LAYER M3 ;
        RECT 10.88 4.836 10.912 10.368 ;
  LAYER M3 ;
        RECT 10.816 4.836 10.848 10.368 ;
  LAYER M3 ;
        RECT 10.752 4.836 10.784 10.368 ;
  LAYER M3 ;
        RECT 10.688 4.836 10.72 10.368 ;
  LAYER M3 ;
        RECT 10.624 4.836 10.656 10.368 ;
  LAYER M3 ;
        RECT 10.56 4.836 10.592 10.368 ;
  LAYER M3 ;
        RECT 10.496 4.836 10.528 10.368 ;
  LAYER M3 ;
        RECT 10.432 4.836 10.464 10.368 ;
  LAYER M3 ;
        RECT 10.368 4.836 10.4 10.368 ;
  LAYER M3 ;
        RECT 10.3 4.836 10.34 10.368 ;
  LAYER M2 ;
        RECT 10.044 10.316 16.036 10.348 ;
  LAYER M2 ;
        RECT 10.044 4.856 16.036 4.888 ;
  LAYER M1 ;
        RECT 21.824 4.836 21.856 10.368 ;
  LAYER M1 ;
        RECT 21.76 4.836 21.792 10.368 ;
  LAYER M1 ;
        RECT 21.696 4.836 21.728 10.368 ;
  LAYER M1 ;
        RECT 21.632 4.836 21.664 10.368 ;
  LAYER M1 ;
        RECT 21.568 4.836 21.6 10.368 ;
  LAYER M1 ;
        RECT 21.504 4.836 21.536 10.368 ;
  LAYER M1 ;
        RECT 21.44 4.836 21.472 10.368 ;
  LAYER M1 ;
        RECT 21.376 4.836 21.408 10.368 ;
  LAYER M1 ;
        RECT 21.312 4.836 21.344 10.368 ;
  LAYER M1 ;
        RECT 21.248 4.836 21.28 10.368 ;
  LAYER M1 ;
        RECT 21.184 4.836 21.216 10.368 ;
  LAYER M1 ;
        RECT 21.12 4.836 21.152 10.368 ;
  LAYER M1 ;
        RECT 21.056 4.836 21.088 10.368 ;
  LAYER M1 ;
        RECT 20.992 4.836 21.024 10.368 ;
  LAYER M1 ;
        RECT 20.928 4.836 20.96 10.368 ;
  LAYER M1 ;
        RECT 20.864 4.836 20.896 10.368 ;
  LAYER M1 ;
        RECT 20.8 4.836 20.832 10.368 ;
  LAYER M1 ;
        RECT 20.736 4.836 20.768 10.368 ;
  LAYER M1 ;
        RECT 20.672 4.836 20.704 10.368 ;
  LAYER M1 ;
        RECT 20.608 4.836 20.64 10.368 ;
  LAYER M1 ;
        RECT 20.544 4.836 20.576 10.368 ;
  LAYER M1 ;
        RECT 20.48 4.836 20.512 10.368 ;
  LAYER M1 ;
        RECT 20.416 4.836 20.448 10.368 ;
  LAYER M1 ;
        RECT 20.352 4.836 20.384 10.368 ;
  LAYER M1 ;
        RECT 20.288 4.836 20.32 10.368 ;
  LAYER M1 ;
        RECT 20.224 4.836 20.256 10.368 ;
  LAYER M1 ;
        RECT 20.16 4.836 20.192 10.368 ;
  LAYER M1 ;
        RECT 20.096 4.836 20.128 10.368 ;
  LAYER M1 ;
        RECT 20.032 4.836 20.064 10.368 ;
  LAYER M1 ;
        RECT 19.968 4.836 20 10.368 ;
  LAYER M1 ;
        RECT 19.904 4.836 19.936 10.368 ;
  LAYER M1 ;
        RECT 19.84 4.836 19.872 10.368 ;
  LAYER M1 ;
        RECT 19.776 4.836 19.808 10.368 ;
  LAYER M1 ;
        RECT 19.712 4.836 19.744 10.368 ;
  LAYER M1 ;
        RECT 19.648 4.836 19.68 10.368 ;
  LAYER M1 ;
        RECT 19.584 4.836 19.616 10.368 ;
  LAYER M1 ;
        RECT 19.52 4.836 19.552 10.368 ;
  LAYER M1 ;
        RECT 19.456 4.836 19.488 10.368 ;
  LAYER M1 ;
        RECT 19.392 4.836 19.424 10.368 ;
  LAYER M1 ;
        RECT 19.328 4.836 19.36 10.368 ;
  LAYER M1 ;
        RECT 19.264 4.836 19.296 10.368 ;
  LAYER M1 ;
        RECT 19.2 4.836 19.232 10.368 ;
  LAYER M1 ;
        RECT 19.136 4.836 19.168 10.368 ;
  LAYER M1 ;
        RECT 19.072 4.836 19.104 10.368 ;
  LAYER M1 ;
        RECT 19.008 4.836 19.04 10.368 ;
  LAYER M1 ;
        RECT 18.944 4.836 18.976 10.368 ;
  LAYER M1 ;
        RECT 18.88 4.836 18.912 10.368 ;
  LAYER M1 ;
        RECT 18.816 4.836 18.848 10.368 ;
  LAYER M1 ;
        RECT 18.752 4.836 18.784 10.368 ;
  LAYER M1 ;
        RECT 18.688 4.836 18.72 10.368 ;
  LAYER M1 ;
        RECT 18.624 4.836 18.656 10.368 ;
  LAYER M1 ;
        RECT 18.56 4.836 18.592 10.368 ;
  LAYER M1 ;
        RECT 18.496 4.836 18.528 10.368 ;
  LAYER M1 ;
        RECT 18.432 4.836 18.464 10.368 ;
  LAYER M1 ;
        RECT 18.368 4.836 18.4 10.368 ;
  LAYER M1 ;
        RECT 18.304 4.836 18.336 10.368 ;
  LAYER M1 ;
        RECT 18.24 4.836 18.272 10.368 ;
  LAYER M1 ;
        RECT 18.176 4.836 18.208 10.368 ;
  LAYER M1 ;
        RECT 18.112 4.836 18.144 10.368 ;
  LAYER M1 ;
        RECT 18.048 4.836 18.08 10.368 ;
  LAYER M1 ;
        RECT 17.984 4.836 18.016 10.368 ;
  LAYER M1 ;
        RECT 17.92 4.836 17.952 10.368 ;
  LAYER M1 ;
        RECT 17.856 4.836 17.888 10.368 ;
  LAYER M1 ;
        RECT 17.792 4.836 17.824 10.368 ;
  LAYER M1 ;
        RECT 17.728 4.836 17.76 10.368 ;
  LAYER M1 ;
        RECT 17.664 4.836 17.696 10.368 ;
  LAYER M1 ;
        RECT 17.6 4.836 17.632 10.368 ;
  LAYER M1 ;
        RECT 17.536 4.836 17.568 10.368 ;
  LAYER M1 ;
        RECT 17.472 4.836 17.504 10.368 ;
  LAYER M1 ;
        RECT 17.408 4.836 17.44 10.368 ;
  LAYER M1 ;
        RECT 17.344 4.836 17.376 10.368 ;
  LAYER M1 ;
        RECT 17.28 4.836 17.312 10.368 ;
  LAYER M1 ;
        RECT 17.216 4.836 17.248 10.368 ;
  LAYER M1 ;
        RECT 17.152 4.836 17.184 10.368 ;
  LAYER M1 ;
        RECT 17.088 4.836 17.12 10.368 ;
  LAYER M1 ;
        RECT 17.024 4.836 17.056 10.368 ;
  LAYER M1 ;
        RECT 16.96 4.836 16.992 10.368 ;
  LAYER M1 ;
        RECT 16.896 4.836 16.928 10.368 ;
  LAYER M1 ;
        RECT 16.832 4.836 16.864 10.368 ;
  LAYER M1 ;
        RECT 16.768 4.836 16.8 10.368 ;
  LAYER M1 ;
        RECT 16.704 4.836 16.736 10.368 ;
  LAYER M1 ;
        RECT 16.64 4.836 16.672 10.368 ;
  LAYER M1 ;
        RECT 16.576 4.836 16.608 10.368 ;
  LAYER M1 ;
        RECT 16.512 4.836 16.544 10.368 ;
  LAYER M1 ;
        RECT 16.448 4.836 16.48 10.368 ;
  LAYER M1 ;
        RECT 16.384 4.836 16.416 10.368 ;
  LAYER M2 ;
        RECT 16.364 4.92 21.876 4.952 ;
  LAYER M2 ;
        RECT 16.364 4.984 21.876 5.016 ;
  LAYER M2 ;
        RECT 16.364 5.048 21.876 5.08 ;
  LAYER M2 ;
        RECT 16.364 5.112 21.876 5.144 ;
  LAYER M2 ;
        RECT 16.364 5.176 21.876 5.208 ;
  LAYER M2 ;
        RECT 16.364 5.24 21.876 5.272 ;
  LAYER M2 ;
        RECT 16.364 5.304 21.876 5.336 ;
  LAYER M2 ;
        RECT 16.364 5.368 21.876 5.4 ;
  LAYER M2 ;
        RECT 16.364 5.432 21.876 5.464 ;
  LAYER M2 ;
        RECT 16.364 5.496 21.876 5.528 ;
  LAYER M2 ;
        RECT 16.364 5.56 21.876 5.592 ;
  LAYER M2 ;
        RECT 16.364 5.624 21.876 5.656 ;
  LAYER M2 ;
        RECT 16.364 5.688 21.876 5.72 ;
  LAYER M2 ;
        RECT 16.364 5.752 21.876 5.784 ;
  LAYER M2 ;
        RECT 16.364 5.816 21.876 5.848 ;
  LAYER M2 ;
        RECT 16.364 5.88 21.876 5.912 ;
  LAYER M2 ;
        RECT 16.364 5.944 21.876 5.976 ;
  LAYER M2 ;
        RECT 16.364 6.008 21.876 6.04 ;
  LAYER M2 ;
        RECT 16.364 6.072 21.876 6.104 ;
  LAYER M2 ;
        RECT 16.364 6.136 21.876 6.168 ;
  LAYER M2 ;
        RECT 16.364 6.2 21.876 6.232 ;
  LAYER M2 ;
        RECT 16.364 6.264 21.876 6.296 ;
  LAYER M2 ;
        RECT 16.364 6.328 21.876 6.36 ;
  LAYER M2 ;
        RECT 16.364 6.392 21.876 6.424 ;
  LAYER M2 ;
        RECT 16.364 6.456 21.876 6.488 ;
  LAYER M2 ;
        RECT 16.364 6.52 21.876 6.552 ;
  LAYER M2 ;
        RECT 16.364 6.584 21.876 6.616 ;
  LAYER M2 ;
        RECT 16.364 6.648 21.876 6.68 ;
  LAYER M2 ;
        RECT 16.364 6.712 21.876 6.744 ;
  LAYER M2 ;
        RECT 16.364 6.776 21.876 6.808 ;
  LAYER M2 ;
        RECT 16.364 6.84 21.876 6.872 ;
  LAYER M2 ;
        RECT 16.364 6.904 21.876 6.936 ;
  LAYER M2 ;
        RECT 16.364 6.968 21.876 7 ;
  LAYER M2 ;
        RECT 16.364 7.032 21.876 7.064 ;
  LAYER M2 ;
        RECT 16.364 7.096 21.876 7.128 ;
  LAYER M2 ;
        RECT 16.364 7.16 21.876 7.192 ;
  LAYER M2 ;
        RECT 16.364 7.224 21.876 7.256 ;
  LAYER M2 ;
        RECT 16.364 7.288 21.876 7.32 ;
  LAYER M2 ;
        RECT 16.364 7.352 21.876 7.384 ;
  LAYER M2 ;
        RECT 16.364 7.416 21.876 7.448 ;
  LAYER M2 ;
        RECT 16.364 7.48 21.876 7.512 ;
  LAYER M2 ;
        RECT 16.364 7.544 21.876 7.576 ;
  LAYER M2 ;
        RECT 16.364 7.608 21.876 7.64 ;
  LAYER M2 ;
        RECT 16.364 7.672 21.876 7.704 ;
  LAYER M2 ;
        RECT 16.364 7.736 21.876 7.768 ;
  LAYER M2 ;
        RECT 16.364 7.8 21.876 7.832 ;
  LAYER M2 ;
        RECT 16.364 7.864 21.876 7.896 ;
  LAYER M2 ;
        RECT 16.364 7.928 21.876 7.96 ;
  LAYER M2 ;
        RECT 16.364 7.992 21.876 8.024 ;
  LAYER M2 ;
        RECT 16.364 8.056 21.876 8.088 ;
  LAYER M2 ;
        RECT 16.364 8.12 21.876 8.152 ;
  LAYER M2 ;
        RECT 16.364 8.184 21.876 8.216 ;
  LAYER M2 ;
        RECT 16.364 8.248 21.876 8.28 ;
  LAYER M2 ;
        RECT 16.364 8.312 21.876 8.344 ;
  LAYER M2 ;
        RECT 16.364 8.376 21.876 8.408 ;
  LAYER M2 ;
        RECT 16.364 8.44 21.876 8.472 ;
  LAYER M2 ;
        RECT 16.364 8.504 21.876 8.536 ;
  LAYER M2 ;
        RECT 16.364 8.568 21.876 8.6 ;
  LAYER M2 ;
        RECT 16.364 8.632 21.876 8.664 ;
  LAYER M2 ;
        RECT 16.364 8.696 21.876 8.728 ;
  LAYER M2 ;
        RECT 16.364 8.76 21.876 8.792 ;
  LAYER M2 ;
        RECT 16.364 8.824 21.876 8.856 ;
  LAYER M2 ;
        RECT 16.364 8.888 21.876 8.92 ;
  LAYER M2 ;
        RECT 16.364 8.952 21.876 8.984 ;
  LAYER M2 ;
        RECT 16.364 9.016 21.876 9.048 ;
  LAYER M2 ;
        RECT 16.364 9.08 21.876 9.112 ;
  LAYER M2 ;
        RECT 16.364 9.144 21.876 9.176 ;
  LAYER M2 ;
        RECT 16.364 9.208 21.876 9.24 ;
  LAYER M2 ;
        RECT 16.364 9.272 21.876 9.304 ;
  LAYER M2 ;
        RECT 16.364 9.336 21.876 9.368 ;
  LAYER M2 ;
        RECT 16.364 9.4 21.876 9.432 ;
  LAYER M2 ;
        RECT 16.364 9.464 21.876 9.496 ;
  LAYER M2 ;
        RECT 16.364 9.528 21.876 9.56 ;
  LAYER M2 ;
        RECT 16.364 9.592 21.876 9.624 ;
  LAYER M2 ;
        RECT 16.364 9.656 21.876 9.688 ;
  LAYER M2 ;
        RECT 16.364 9.72 21.876 9.752 ;
  LAYER M2 ;
        RECT 16.364 9.784 21.876 9.816 ;
  LAYER M2 ;
        RECT 16.364 9.848 21.876 9.88 ;
  LAYER M2 ;
        RECT 16.364 9.912 21.876 9.944 ;
  LAYER M2 ;
        RECT 16.364 9.976 21.876 10.008 ;
  LAYER M2 ;
        RECT 16.364 10.04 21.876 10.072 ;
  LAYER M2 ;
        RECT 16.364 10.104 21.876 10.136 ;
  LAYER M2 ;
        RECT 16.364 10.168 21.876 10.2 ;
  LAYER M2 ;
        RECT 16.364 10.232 21.876 10.264 ;
  LAYER M3 ;
        RECT 21.824 4.836 21.856 10.368 ;
  LAYER M3 ;
        RECT 21.76 4.836 21.792 10.368 ;
  LAYER M3 ;
        RECT 21.696 4.836 21.728 10.368 ;
  LAYER M3 ;
        RECT 21.632 4.836 21.664 10.368 ;
  LAYER M3 ;
        RECT 21.568 4.836 21.6 10.368 ;
  LAYER M3 ;
        RECT 21.504 4.836 21.536 10.368 ;
  LAYER M3 ;
        RECT 21.44 4.836 21.472 10.368 ;
  LAYER M3 ;
        RECT 21.376 4.836 21.408 10.368 ;
  LAYER M3 ;
        RECT 21.312 4.836 21.344 10.368 ;
  LAYER M3 ;
        RECT 21.248 4.836 21.28 10.368 ;
  LAYER M3 ;
        RECT 21.184 4.836 21.216 10.368 ;
  LAYER M3 ;
        RECT 21.12 4.836 21.152 10.368 ;
  LAYER M3 ;
        RECT 21.056 4.836 21.088 10.368 ;
  LAYER M3 ;
        RECT 20.992 4.836 21.024 10.368 ;
  LAYER M3 ;
        RECT 20.928 4.836 20.96 10.368 ;
  LAYER M3 ;
        RECT 20.864 4.836 20.896 10.368 ;
  LAYER M3 ;
        RECT 20.8 4.836 20.832 10.368 ;
  LAYER M3 ;
        RECT 20.736 4.836 20.768 10.368 ;
  LAYER M3 ;
        RECT 20.672 4.836 20.704 10.368 ;
  LAYER M3 ;
        RECT 20.608 4.836 20.64 10.368 ;
  LAYER M3 ;
        RECT 20.544 4.836 20.576 10.368 ;
  LAYER M3 ;
        RECT 20.48 4.836 20.512 10.368 ;
  LAYER M3 ;
        RECT 20.416 4.836 20.448 10.368 ;
  LAYER M3 ;
        RECT 20.352 4.836 20.384 10.368 ;
  LAYER M3 ;
        RECT 20.288 4.836 20.32 10.368 ;
  LAYER M3 ;
        RECT 20.224 4.836 20.256 10.368 ;
  LAYER M3 ;
        RECT 20.16 4.836 20.192 10.368 ;
  LAYER M3 ;
        RECT 20.096 4.836 20.128 10.368 ;
  LAYER M3 ;
        RECT 20.032 4.836 20.064 10.368 ;
  LAYER M3 ;
        RECT 19.968 4.836 20 10.368 ;
  LAYER M3 ;
        RECT 19.904 4.836 19.936 10.368 ;
  LAYER M3 ;
        RECT 19.84 4.836 19.872 10.368 ;
  LAYER M3 ;
        RECT 19.776 4.836 19.808 10.368 ;
  LAYER M3 ;
        RECT 19.712 4.836 19.744 10.368 ;
  LAYER M3 ;
        RECT 19.648 4.836 19.68 10.368 ;
  LAYER M3 ;
        RECT 19.584 4.836 19.616 10.368 ;
  LAYER M3 ;
        RECT 19.52 4.836 19.552 10.368 ;
  LAYER M3 ;
        RECT 19.456 4.836 19.488 10.368 ;
  LAYER M3 ;
        RECT 19.392 4.836 19.424 10.368 ;
  LAYER M3 ;
        RECT 19.328 4.836 19.36 10.368 ;
  LAYER M3 ;
        RECT 19.264 4.836 19.296 10.368 ;
  LAYER M3 ;
        RECT 19.2 4.836 19.232 10.368 ;
  LAYER M3 ;
        RECT 19.136 4.836 19.168 10.368 ;
  LAYER M3 ;
        RECT 19.072 4.836 19.104 10.368 ;
  LAYER M3 ;
        RECT 19.008 4.836 19.04 10.368 ;
  LAYER M3 ;
        RECT 18.944 4.836 18.976 10.368 ;
  LAYER M3 ;
        RECT 18.88 4.836 18.912 10.368 ;
  LAYER M3 ;
        RECT 18.816 4.836 18.848 10.368 ;
  LAYER M3 ;
        RECT 18.752 4.836 18.784 10.368 ;
  LAYER M3 ;
        RECT 18.688 4.836 18.72 10.368 ;
  LAYER M3 ;
        RECT 18.624 4.836 18.656 10.368 ;
  LAYER M3 ;
        RECT 18.56 4.836 18.592 10.368 ;
  LAYER M3 ;
        RECT 18.496 4.836 18.528 10.368 ;
  LAYER M3 ;
        RECT 18.432 4.836 18.464 10.368 ;
  LAYER M3 ;
        RECT 18.368 4.836 18.4 10.368 ;
  LAYER M3 ;
        RECT 18.304 4.836 18.336 10.368 ;
  LAYER M3 ;
        RECT 18.24 4.836 18.272 10.368 ;
  LAYER M3 ;
        RECT 18.176 4.836 18.208 10.368 ;
  LAYER M3 ;
        RECT 18.112 4.836 18.144 10.368 ;
  LAYER M3 ;
        RECT 18.048 4.836 18.08 10.368 ;
  LAYER M3 ;
        RECT 17.984 4.836 18.016 10.368 ;
  LAYER M3 ;
        RECT 17.92 4.836 17.952 10.368 ;
  LAYER M3 ;
        RECT 17.856 4.836 17.888 10.368 ;
  LAYER M3 ;
        RECT 17.792 4.836 17.824 10.368 ;
  LAYER M3 ;
        RECT 17.728 4.836 17.76 10.368 ;
  LAYER M3 ;
        RECT 17.664 4.836 17.696 10.368 ;
  LAYER M3 ;
        RECT 17.6 4.836 17.632 10.368 ;
  LAYER M3 ;
        RECT 17.536 4.836 17.568 10.368 ;
  LAYER M3 ;
        RECT 17.472 4.836 17.504 10.368 ;
  LAYER M3 ;
        RECT 17.408 4.836 17.44 10.368 ;
  LAYER M3 ;
        RECT 17.344 4.836 17.376 10.368 ;
  LAYER M3 ;
        RECT 17.28 4.836 17.312 10.368 ;
  LAYER M3 ;
        RECT 17.216 4.836 17.248 10.368 ;
  LAYER M3 ;
        RECT 17.152 4.836 17.184 10.368 ;
  LAYER M3 ;
        RECT 17.088 4.836 17.12 10.368 ;
  LAYER M3 ;
        RECT 17.024 4.836 17.056 10.368 ;
  LAYER M3 ;
        RECT 16.96 4.836 16.992 10.368 ;
  LAYER M3 ;
        RECT 16.896 4.836 16.928 10.368 ;
  LAYER M3 ;
        RECT 16.832 4.836 16.864 10.368 ;
  LAYER M3 ;
        RECT 16.768 4.836 16.8 10.368 ;
  LAYER M3 ;
        RECT 16.704 4.836 16.736 10.368 ;
  LAYER M3 ;
        RECT 16.64 4.836 16.672 10.368 ;
  LAYER M3 ;
        RECT 16.576 4.836 16.608 10.368 ;
  LAYER M3 ;
        RECT 16.512 4.836 16.544 10.368 ;
  LAYER M3 ;
        RECT 16.448 4.836 16.48 10.368 ;
  LAYER M3 ;
        RECT 16.38 4.836 16.42 10.368 ;
  LAYER M2 ;
        RECT 16.124 10.316 22.116 10.348 ;
  LAYER M2 ;
        RECT 16.124 4.856 22.116 4.888 ;
  LAYER M1 ;
        RECT 36.064 4.836 36.096 10.368 ;
  LAYER M1 ;
        RECT 36 4.836 36.032 10.368 ;
  LAYER M1 ;
        RECT 35.936 4.836 35.968 10.368 ;
  LAYER M1 ;
        RECT 35.872 4.836 35.904 10.368 ;
  LAYER M1 ;
        RECT 35.808 4.836 35.84 10.368 ;
  LAYER M1 ;
        RECT 35.744 4.836 35.776 10.368 ;
  LAYER M1 ;
        RECT 35.68 4.836 35.712 10.368 ;
  LAYER M1 ;
        RECT 35.616 4.836 35.648 10.368 ;
  LAYER M1 ;
        RECT 35.552 4.836 35.584 10.368 ;
  LAYER M1 ;
        RECT 35.488 4.836 35.52 10.368 ;
  LAYER M1 ;
        RECT 35.424 4.836 35.456 10.368 ;
  LAYER M1 ;
        RECT 35.36 4.836 35.392 10.368 ;
  LAYER M1 ;
        RECT 35.296 4.836 35.328 10.368 ;
  LAYER M1 ;
        RECT 35.232 4.836 35.264 10.368 ;
  LAYER M1 ;
        RECT 35.168 4.836 35.2 10.368 ;
  LAYER M1 ;
        RECT 35.104 4.836 35.136 10.368 ;
  LAYER M1 ;
        RECT 35.04 4.836 35.072 10.368 ;
  LAYER M1 ;
        RECT 34.976 4.836 35.008 10.368 ;
  LAYER M1 ;
        RECT 34.912 4.836 34.944 10.368 ;
  LAYER M1 ;
        RECT 34.848 4.836 34.88 10.368 ;
  LAYER M1 ;
        RECT 34.784 4.836 34.816 10.368 ;
  LAYER M1 ;
        RECT 34.72 4.836 34.752 10.368 ;
  LAYER M1 ;
        RECT 34.656 4.836 34.688 10.368 ;
  LAYER M1 ;
        RECT 34.592 4.836 34.624 10.368 ;
  LAYER M1 ;
        RECT 34.528 4.836 34.56 10.368 ;
  LAYER M1 ;
        RECT 34.464 4.836 34.496 10.368 ;
  LAYER M1 ;
        RECT 34.4 4.836 34.432 10.368 ;
  LAYER M1 ;
        RECT 34.336 4.836 34.368 10.368 ;
  LAYER M1 ;
        RECT 34.272 4.836 34.304 10.368 ;
  LAYER M1 ;
        RECT 34.208 4.836 34.24 10.368 ;
  LAYER M1 ;
        RECT 34.144 4.836 34.176 10.368 ;
  LAYER M1 ;
        RECT 34.08 4.836 34.112 10.368 ;
  LAYER M1 ;
        RECT 34.016 4.836 34.048 10.368 ;
  LAYER M1 ;
        RECT 33.952 4.836 33.984 10.368 ;
  LAYER M1 ;
        RECT 33.888 4.836 33.92 10.368 ;
  LAYER M1 ;
        RECT 33.824 4.836 33.856 10.368 ;
  LAYER M1 ;
        RECT 33.76 4.836 33.792 10.368 ;
  LAYER M1 ;
        RECT 33.696 4.836 33.728 10.368 ;
  LAYER M1 ;
        RECT 33.632 4.836 33.664 10.368 ;
  LAYER M1 ;
        RECT 33.568 4.836 33.6 10.368 ;
  LAYER M1 ;
        RECT 33.504 4.836 33.536 10.368 ;
  LAYER M1 ;
        RECT 33.44 4.836 33.472 10.368 ;
  LAYER M1 ;
        RECT 33.376 4.836 33.408 10.368 ;
  LAYER M1 ;
        RECT 33.312 4.836 33.344 10.368 ;
  LAYER M1 ;
        RECT 33.248 4.836 33.28 10.368 ;
  LAYER M1 ;
        RECT 33.184 4.836 33.216 10.368 ;
  LAYER M1 ;
        RECT 33.12 4.836 33.152 10.368 ;
  LAYER M1 ;
        RECT 33.056 4.836 33.088 10.368 ;
  LAYER M1 ;
        RECT 32.992 4.836 33.024 10.368 ;
  LAYER M1 ;
        RECT 32.928 4.836 32.96 10.368 ;
  LAYER M1 ;
        RECT 32.864 4.836 32.896 10.368 ;
  LAYER M1 ;
        RECT 32.8 4.836 32.832 10.368 ;
  LAYER M1 ;
        RECT 32.736 4.836 32.768 10.368 ;
  LAYER M1 ;
        RECT 32.672 4.836 32.704 10.368 ;
  LAYER M1 ;
        RECT 32.608 4.836 32.64 10.368 ;
  LAYER M1 ;
        RECT 32.544 4.836 32.576 10.368 ;
  LAYER M1 ;
        RECT 32.48 4.836 32.512 10.368 ;
  LAYER M1 ;
        RECT 32.416 4.836 32.448 10.368 ;
  LAYER M1 ;
        RECT 32.352 4.836 32.384 10.368 ;
  LAYER M1 ;
        RECT 32.288 4.836 32.32 10.368 ;
  LAYER M1 ;
        RECT 32.224 4.836 32.256 10.368 ;
  LAYER M1 ;
        RECT 32.16 4.836 32.192 10.368 ;
  LAYER M1 ;
        RECT 32.096 4.836 32.128 10.368 ;
  LAYER M1 ;
        RECT 32.032 4.836 32.064 10.368 ;
  LAYER M1 ;
        RECT 31.968 4.836 32 10.368 ;
  LAYER M1 ;
        RECT 31.904 4.836 31.936 10.368 ;
  LAYER M1 ;
        RECT 31.84 4.836 31.872 10.368 ;
  LAYER M1 ;
        RECT 31.776 4.836 31.808 10.368 ;
  LAYER M1 ;
        RECT 31.712 4.836 31.744 10.368 ;
  LAYER M1 ;
        RECT 31.648 4.836 31.68 10.368 ;
  LAYER M1 ;
        RECT 31.584 4.836 31.616 10.368 ;
  LAYER M1 ;
        RECT 31.52 4.836 31.552 10.368 ;
  LAYER M1 ;
        RECT 31.456 4.836 31.488 10.368 ;
  LAYER M1 ;
        RECT 31.392 4.836 31.424 10.368 ;
  LAYER M1 ;
        RECT 31.328 4.836 31.36 10.368 ;
  LAYER M1 ;
        RECT 31.264 4.836 31.296 10.368 ;
  LAYER M1 ;
        RECT 31.2 4.836 31.232 10.368 ;
  LAYER M1 ;
        RECT 31.136 4.836 31.168 10.368 ;
  LAYER M1 ;
        RECT 31.072 4.836 31.104 10.368 ;
  LAYER M1 ;
        RECT 31.008 4.836 31.04 10.368 ;
  LAYER M1 ;
        RECT 30.944 4.836 30.976 10.368 ;
  LAYER M1 ;
        RECT 30.88 4.836 30.912 10.368 ;
  LAYER M1 ;
        RECT 30.816 4.836 30.848 10.368 ;
  LAYER M1 ;
        RECT 30.752 4.836 30.784 10.368 ;
  LAYER M1 ;
        RECT 30.688 4.836 30.72 10.368 ;
  LAYER M1 ;
        RECT 30.624 4.836 30.656 10.368 ;
  LAYER M2 ;
        RECT 30.604 10.252 36.116 10.284 ;
  LAYER M2 ;
        RECT 30.604 10.188 36.116 10.22 ;
  LAYER M2 ;
        RECT 30.604 10.124 36.116 10.156 ;
  LAYER M2 ;
        RECT 30.604 10.06 36.116 10.092 ;
  LAYER M2 ;
        RECT 30.604 9.996 36.116 10.028 ;
  LAYER M2 ;
        RECT 30.604 9.932 36.116 9.964 ;
  LAYER M2 ;
        RECT 30.604 9.868 36.116 9.9 ;
  LAYER M2 ;
        RECT 30.604 9.804 36.116 9.836 ;
  LAYER M2 ;
        RECT 30.604 9.74 36.116 9.772 ;
  LAYER M2 ;
        RECT 30.604 9.676 36.116 9.708 ;
  LAYER M2 ;
        RECT 30.604 9.612 36.116 9.644 ;
  LAYER M2 ;
        RECT 30.604 9.548 36.116 9.58 ;
  LAYER M2 ;
        RECT 30.604 9.484 36.116 9.516 ;
  LAYER M2 ;
        RECT 30.604 9.42 36.116 9.452 ;
  LAYER M2 ;
        RECT 30.604 9.356 36.116 9.388 ;
  LAYER M2 ;
        RECT 30.604 9.292 36.116 9.324 ;
  LAYER M2 ;
        RECT 30.604 9.228 36.116 9.26 ;
  LAYER M2 ;
        RECT 30.604 9.164 36.116 9.196 ;
  LAYER M2 ;
        RECT 30.604 9.1 36.116 9.132 ;
  LAYER M2 ;
        RECT 30.604 9.036 36.116 9.068 ;
  LAYER M2 ;
        RECT 30.604 8.972 36.116 9.004 ;
  LAYER M2 ;
        RECT 30.604 8.908 36.116 8.94 ;
  LAYER M2 ;
        RECT 30.604 8.844 36.116 8.876 ;
  LAYER M2 ;
        RECT 30.604 8.78 36.116 8.812 ;
  LAYER M2 ;
        RECT 30.604 8.716 36.116 8.748 ;
  LAYER M2 ;
        RECT 30.604 8.652 36.116 8.684 ;
  LAYER M2 ;
        RECT 30.604 8.588 36.116 8.62 ;
  LAYER M2 ;
        RECT 30.604 8.524 36.116 8.556 ;
  LAYER M2 ;
        RECT 30.604 8.46 36.116 8.492 ;
  LAYER M2 ;
        RECT 30.604 8.396 36.116 8.428 ;
  LAYER M2 ;
        RECT 30.604 8.332 36.116 8.364 ;
  LAYER M2 ;
        RECT 30.604 8.268 36.116 8.3 ;
  LAYER M2 ;
        RECT 30.604 8.204 36.116 8.236 ;
  LAYER M2 ;
        RECT 30.604 8.14 36.116 8.172 ;
  LAYER M2 ;
        RECT 30.604 8.076 36.116 8.108 ;
  LAYER M2 ;
        RECT 30.604 8.012 36.116 8.044 ;
  LAYER M2 ;
        RECT 30.604 7.948 36.116 7.98 ;
  LAYER M2 ;
        RECT 30.604 7.884 36.116 7.916 ;
  LAYER M2 ;
        RECT 30.604 7.82 36.116 7.852 ;
  LAYER M2 ;
        RECT 30.604 7.756 36.116 7.788 ;
  LAYER M2 ;
        RECT 30.604 7.692 36.116 7.724 ;
  LAYER M2 ;
        RECT 30.604 7.628 36.116 7.66 ;
  LAYER M2 ;
        RECT 30.604 7.564 36.116 7.596 ;
  LAYER M2 ;
        RECT 30.604 7.5 36.116 7.532 ;
  LAYER M2 ;
        RECT 30.604 7.436 36.116 7.468 ;
  LAYER M2 ;
        RECT 30.604 7.372 36.116 7.404 ;
  LAYER M2 ;
        RECT 30.604 7.308 36.116 7.34 ;
  LAYER M2 ;
        RECT 30.604 7.244 36.116 7.276 ;
  LAYER M2 ;
        RECT 30.604 7.18 36.116 7.212 ;
  LAYER M2 ;
        RECT 30.604 7.116 36.116 7.148 ;
  LAYER M2 ;
        RECT 30.604 7.052 36.116 7.084 ;
  LAYER M2 ;
        RECT 30.604 6.988 36.116 7.02 ;
  LAYER M2 ;
        RECT 30.604 6.924 36.116 6.956 ;
  LAYER M2 ;
        RECT 30.604 6.86 36.116 6.892 ;
  LAYER M2 ;
        RECT 30.604 6.796 36.116 6.828 ;
  LAYER M2 ;
        RECT 30.604 6.732 36.116 6.764 ;
  LAYER M2 ;
        RECT 30.604 6.668 36.116 6.7 ;
  LAYER M2 ;
        RECT 30.604 6.604 36.116 6.636 ;
  LAYER M2 ;
        RECT 30.604 6.54 36.116 6.572 ;
  LAYER M2 ;
        RECT 30.604 6.476 36.116 6.508 ;
  LAYER M2 ;
        RECT 30.604 6.412 36.116 6.444 ;
  LAYER M2 ;
        RECT 30.604 6.348 36.116 6.38 ;
  LAYER M2 ;
        RECT 30.604 6.284 36.116 6.316 ;
  LAYER M2 ;
        RECT 30.604 6.22 36.116 6.252 ;
  LAYER M2 ;
        RECT 30.604 6.156 36.116 6.188 ;
  LAYER M2 ;
        RECT 30.604 6.092 36.116 6.124 ;
  LAYER M2 ;
        RECT 30.604 6.028 36.116 6.06 ;
  LAYER M2 ;
        RECT 30.604 5.964 36.116 5.996 ;
  LAYER M2 ;
        RECT 30.604 5.9 36.116 5.932 ;
  LAYER M2 ;
        RECT 30.604 5.836 36.116 5.868 ;
  LAYER M2 ;
        RECT 30.604 5.772 36.116 5.804 ;
  LAYER M2 ;
        RECT 30.604 5.708 36.116 5.74 ;
  LAYER M2 ;
        RECT 30.604 5.644 36.116 5.676 ;
  LAYER M2 ;
        RECT 30.604 5.58 36.116 5.612 ;
  LAYER M2 ;
        RECT 30.604 5.516 36.116 5.548 ;
  LAYER M2 ;
        RECT 30.604 5.452 36.116 5.484 ;
  LAYER M2 ;
        RECT 30.604 5.388 36.116 5.42 ;
  LAYER M2 ;
        RECT 30.604 5.324 36.116 5.356 ;
  LAYER M2 ;
        RECT 30.604 5.26 36.116 5.292 ;
  LAYER M2 ;
        RECT 30.604 5.196 36.116 5.228 ;
  LAYER M2 ;
        RECT 30.604 5.132 36.116 5.164 ;
  LAYER M2 ;
        RECT 30.604 5.068 36.116 5.1 ;
  LAYER M2 ;
        RECT 30.604 5.004 36.116 5.036 ;
  LAYER M2 ;
        RECT 30.604 4.94 36.116 4.972 ;
  LAYER M3 ;
        RECT 36.064 4.836 36.096 10.368 ;
  LAYER M3 ;
        RECT 36 4.836 36.032 10.368 ;
  LAYER M3 ;
        RECT 35.936 4.836 35.968 10.368 ;
  LAYER M3 ;
        RECT 35.872 4.836 35.904 10.368 ;
  LAYER M3 ;
        RECT 35.808 4.836 35.84 10.368 ;
  LAYER M3 ;
        RECT 35.744 4.836 35.776 10.368 ;
  LAYER M3 ;
        RECT 35.68 4.836 35.712 10.368 ;
  LAYER M3 ;
        RECT 35.616 4.836 35.648 10.368 ;
  LAYER M3 ;
        RECT 35.552 4.836 35.584 10.368 ;
  LAYER M3 ;
        RECT 35.488 4.836 35.52 10.368 ;
  LAYER M3 ;
        RECT 35.424 4.836 35.456 10.368 ;
  LAYER M3 ;
        RECT 35.36 4.836 35.392 10.368 ;
  LAYER M3 ;
        RECT 35.296 4.836 35.328 10.368 ;
  LAYER M3 ;
        RECT 35.232 4.836 35.264 10.368 ;
  LAYER M3 ;
        RECT 35.168 4.836 35.2 10.368 ;
  LAYER M3 ;
        RECT 35.104 4.836 35.136 10.368 ;
  LAYER M3 ;
        RECT 35.04 4.836 35.072 10.368 ;
  LAYER M3 ;
        RECT 34.976 4.836 35.008 10.368 ;
  LAYER M3 ;
        RECT 34.912 4.836 34.944 10.368 ;
  LAYER M3 ;
        RECT 34.848 4.836 34.88 10.368 ;
  LAYER M3 ;
        RECT 34.784 4.836 34.816 10.368 ;
  LAYER M3 ;
        RECT 34.72 4.836 34.752 10.368 ;
  LAYER M3 ;
        RECT 34.656 4.836 34.688 10.368 ;
  LAYER M3 ;
        RECT 34.592 4.836 34.624 10.368 ;
  LAYER M3 ;
        RECT 34.528 4.836 34.56 10.368 ;
  LAYER M3 ;
        RECT 34.464 4.836 34.496 10.368 ;
  LAYER M3 ;
        RECT 34.4 4.836 34.432 10.368 ;
  LAYER M3 ;
        RECT 34.336 4.836 34.368 10.368 ;
  LAYER M3 ;
        RECT 34.272 4.836 34.304 10.368 ;
  LAYER M3 ;
        RECT 34.208 4.836 34.24 10.368 ;
  LAYER M3 ;
        RECT 34.144 4.836 34.176 10.368 ;
  LAYER M3 ;
        RECT 34.08 4.836 34.112 10.368 ;
  LAYER M3 ;
        RECT 34.016 4.836 34.048 10.368 ;
  LAYER M3 ;
        RECT 33.952 4.836 33.984 10.368 ;
  LAYER M3 ;
        RECT 33.888 4.836 33.92 10.368 ;
  LAYER M3 ;
        RECT 33.824 4.836 33.856 10.368 ;
  LAYER M3 ;
        RECT 33.76 4.836 33.792 10.368 ;
  LAYER M3 ;
        RECT 33.696 4.836 33.728 10.368 ;
  LAYER M3 ;
        RECT 33.632 4.836 33.664 10.368 ;
  LAYER M3 ;
        RECT 33.568 4.836 33.6 10.368 ;
  LAYER M3 ;
        RECT 33.504 4.836 33.536 10.368 ;
  LAYER M3 ;
        RECT 33.44 4.836 33.472 10.368 ;
  LAYER M3 ;
        RECT 33.376 4.836 33.408 10.368 ;
  LAYER M3 ;
        RECT 33.312 4.836 33.344 10.368 ;
  LAYER M3 ;
        RECT 33.248 4.836 33.28 10.368 ;
  LAYER M3 ;
        RECT 33.184 4.836 33.216 10.368 ;
  LAYER M3 ;
        RECT 33.12 4.836 33.152 10.368 ;
  LAYER M3 ;
        RECT 33.056 4.836 33.088 10.368 ;
  LAYER M3 ;
        RECT 32.992 4.836 33.024 10.368 ;
  LAYER M3 ;
        RECT 32.928 4.836 32.96 10.368 ;
  LAYER M3 ;
        RECT 32.864 4.836 32.896 10.368 ;
  LAYER M3 ;
        RECT 32.8 4.836 32.832 10.368 ;
  LAYER M3 ;
        RECT 32.736 4.836 32.768 10.368 ;
  LAYER M3 ;
        RECT 32.672 4.836 32.704 10.368 ;
  LAYER M3 ;
        RECT 32.608 4.836 32.64 10.368 ;
  LAYER M3 ;
        RECT 32.544 4.836 32.576 10.368 ;
  LAYER M3 ;
        RECT 32.48 4.836 32.512 10.368 ;
  LAYER M3 ;
        RECT 32.416 4.836 32.448 10.368 ;
  LAYER M3 ;
        RECT 32.352 4.836 32.384 10.368 ;
  LAYER M3 ;
        RECT 32.288 4.836 32.32 10.368 ;
  LAYER M3 ;
        RECT 32.224 4.836 32.256 10.368 ;
  LAYER M3 ;
        RECT 32.16 4.836 32.192 10.368 ;
  LAYER M3 ;
        RECT 32.096 4.836 32.128 10.368 ;
  LAYER M3 ;
        RECT 32.032 4.836 32.064 10.368 ;
  LAYER M3 ;
        RECT 31.968 4.836 32 10.368 ;
  LAYER M3 ;
        RECT 31.904 4.836 31.936 10.368 ;
  LAYER M3 ;
        RECT 31.84 4.836 31.872 10.368 ;
  LAYER M3 ;
        RECT 31.776 4.836 31.808 10.368 ;
  LAYER M3 ;
        RECT 31.712 4.836 31.744 10.368 ;
  LAYER M3 ;
        RECT 31.648 4.836 31.68 10.368 ;
  LAYER M3 ;
        RECT 31.584 4.836 31.616 10.368 ;
  LAYER M3 ;
        RECT 31.52 4.836 31.552 10.368 ;
  LAYER M3 ;
        RECT 31.456 4.836 31.488 10.368 ;
  LAYER M3 ;
        RECT 31.392 4.836 31.424 10.368 ;
  LAYER M3 ;
        RECT 31.328 4.836 31.36 10.368 ;
  LAYER M3 ;
        RECT 31.264 4.836 31.296 10.368 ;
  LAYER M3 ;
        RECT 31.2 4.836 31.232 10.368 ;
  LAYER M3 ;
        RECT 31.136 4.836 31.168 10.368 ;
  LAYER M3 ;
        RECT 31.072 4.836 31.104 10.368 ;
  LAYER M3 ;
        RECT 31.008 4.836 31.04 10.368 ;
  LAYER M3 ;
        RECT 30.944 4.836 30.976 10.368 ;
  LAYER M3 ;
        RECT 30.88 4.836 30.912 10.368 ;
  LAYER M3 ;
        RECT 30.816 4.836 30.848 10.368 ;
  LAYER M3 ;
        RECT 30.752 4.836 30.784 10.368 ;
  LAYER M3 ;
        RECT 30.688 4.836 30.72 10.368 ;
  LAYER M3 ;
        RECT 30.62 4.836 30.66 10.368 ;
  LAYER M2 ;
        RECT 30.364 4.856 36.356 4.888 ;
  LAYER M2 ;
        RECT 30.364 10.316 36.356 10.348 ;
  LAYER M1 ;
        RECT 22.464 4.836 22.496 10.368 ;
  LAYER M1 ;
        RECT 22.528 4.836 22.56 10.368 ;
  LAYER M1 ;
        RECT 22.592 4.836 22.624 10.368 ;
  LAYER M1 ;
        RECT 22.656 4.836 22.688 10.368 ;
  LAYER M1 ;
        RECT 22.72 4.836 22.752 10.368 ;
  LAYER M1 ;
        RECT 22.784 4.836 22.816 10.368 ;
  LAYER M1 ;
        RECT 22.848 4.836 22.88 10.368 ;
  LAYER M1 ;
        RECT 22.912 4.836 22.944 10.368 ;
  LAYER M1 ;
        RECT 22.976 4.836 23.008 10.368 ;
  LAYER M1 ;
        RECT 23.04 4.836 23.072 10.368 ;
  LAYER M1 ;
        RECT 23.104 4.836 23.136 10.368 ;
  LAYER M1 ;
        RECT 23.168 4.836 23.2 10.368 ;
  LAYER M1 ;
        RECT 23.232 4.836 23.264 10.368 ;
  LAYER M1 ;
        RECT 23.296 4.836 23.328 10.368 ;
  LAYER M1 ;
        RECT 23.36 4.836 23.392 10.368 ;
  LAYER M1 ;
        RECT 23.424 4.836 23.456 10.368 ;
  LAYER M1 ;
        RECT 23.488 4.836 23.52 10.368 ;
  LAYER M1 ;
        RECT 23.552 4.836 23.584 10.368 ;
  LAYER M1 ;
        RECT 23.616 4.836 23.648 10.368 ;
  LAYER M1 ;
        RECT 23.68 4.836 23.712 10.368 ;
  LAYER M1 ;
        RECT 23.744 4.836 23.776 10.368 ;
  LAYER M1 ;
        RECT 23.808 4.836 23.84 10.368 ;
  LAYER M1 ;
        RECT 23.872 4.836 23.904 10.368 ;
  LAYER M1 ;
        RECT 23.936 4.836 23.968 10.368 ;
  LAYER M1 ;
        RECT 24 4.836 24.032 10.368 ;
  LAYER M1 ;
        RECT 24.064 4.836 24.096 10.368 ;
  LAYER M1 ;
        RECT 24.128 4.836 24.16 10.368 ;
  LAYER M1 ;
        RECT 24.192 4.836 24.224 10.368 ;
  LAYER M1 ;
        RECT 24.256 4.836 24.288 10.368 ;
  LAYER M1 ;
        RECT 24.32 4.836 24.352 10.368 ;
  LAYER M1 ;
        RECT 24.384 4.836 24.416 10.368 ;
  LAYER M1 ;
        RECT 24.448 4.836 24.48 10.368 ;
  LAYER M1 ;
        RECT 24.512 4.836 24.544 10.368 ;
  LAYER M1 ;
        RECT 24.576 4.836 24.608 10.368 ;
  LAYER M1 ;
        RECT 24.64 4.836 24.672 10.368 ;
  LAYER M1 ;
        RECT 24.704 4.836 24.736 10.368 ;
  LAYER M1 ;
        RECT 24.768 4.836 24.8 10.368 ;
  LAYER M1 ;
        RECT 24.832 4.836 24.864 10.368 ;
  LAYER M1 ;
        RECT 24.896 4.836 24.928 10.368 ;
  LAYER M1 ;
        RECT 24.96 4.836 24.992 10.368 ;
  LAYER M1 ;
        RECT 25.024 4.836 25.056 10.368 ;
  LAYER M1 ;
        RECT 25.088 4.836 25.12 10.368 ;
  LAYER M1 ;
        RECT 25.152 4.836 25.184 10.368 ;
  LAYER M1 ;
        RECT 25.216 4.836 25.248 10.368 ;
  LAYER M1 ;
        RECT 25.28 4.836 25.312 10.368 ;
  LAYER M1 ;
        RECT 25.344 4.836 25.376 10.368 ;
  LAYER M1 ;
        RECT 25.408 4.836 25.44 10.368 ;
  LAYER M1 ;
        RECT 25.472 4.836 25.504 10.368 ;
  LAYER M1 ;
        RECT 25.536 4.836 25.568 10.368 ;
  LAYER M1 ;
        RECT 25.6 4.836 25.632 10.368 ;
  LAYER M1 ;
        RECT 25.664 4.836 25.696 10.368 ;
  LAYER M1 ;
        RECT 25.728 4.836 25.76 10.368 ;
  LAYER M1 ;
        RECT 25.792 4.836 25.824 10.368 ;
  LAYER M1 ;
        RECT 25.856 4.836 25.888 10.368 ;
  LAYER M1 ;
        RECT 25.92 4.836 25.952 10.368 ;
  LAYER M1 ;
        RECT 25.984 4.836 26.016 10.368 ;
  LAYER M1 ;
        RECT 26.048 4.836 26.08 10.368 ;
  LAYER M1 ;
        RECT 26.112 4.836 26.144 10.368 ;
  LAYER M1 ;
        RECT 26.176 4.836 26.208 10.368 ;
  LAYER M1 ;
        RECT 26.24 4.836 26.272 10.368 ;
  LAYER M1 ;
        RECT 26.304 4.836 26.336 10.368 ;
  LAYER M1 ;
        RECT 26.368 4.836 26.4 10.368 ;
  LAYER M1 ;
        RECT 26.432 4.836 26.464 10.368 ;
  LAYER M1 ;
        RECT 26.496 4.836 26.528 10.368 ;
  LAYER M1 ;
        RECT 26.56 4.836 26.592 10.368 ;
  LAYER M1 ;
        RECT 26.624 4.836 26.656 10.368 ;
  LAYER M1 ;
        RECT 26.688 4.836 26.72 10.368 ;
  LAYER M1 ;
        RECT 26.752 4.836 26.784 10.368 ;
  LAYER M1 ;
        RECT 26.816 4.836 26.848 10.368 ;
  LAYER M1 ;
        RECT 26.88 4.836 26.912 10.368 ;
  LAYER M1 ;
        RECT 26.944 4.836 26.976 10.368 ;
  LAYER M1 ;
        RECT 27.008 4.836 27.04 10.368 ;
  LAYER M1 ;
        RECT 27.072 4.836 27.104 10.368 ;
  LAYER M1 ;
        RECT 27.136 4.836 27.168 10.368 ;
  LAYER M1 ;
        RECT 27.2 4.836 27.232 10.368 ;
  LAYER M1 ;
        RECT 27.264 4.836 27.296 10.368 ;
  LAYER M1 ;
        RECT 27.328 4.836 27.36 10.368 ;
  LAYER M1 ;
        RECT 27.392 4.836 27.424 10.368 ;
  LAYER M1 ;
        RECT 27.456 4.836 27.488 10.368 ;
  LAYER M1 ;
        RECT 27.52 4.836 27.552 10.368 ;
  LAYER M1 ;
        RECT 27.584 4.836 27.616 10.368 ;
  LAYER M1 ;
        RECT 27.648 4.836 27.68 10.368 ;
  LAYER M1 ;
        RECT 27.712 4.836 27.744 10.368 ;
  LAYER M1 ;
        RECT 27.776 4.836 27.808 10.368 ;
  LAYER M1 ;
        RECT 27.84 4.836 27.872 10.368 ;
  LAYER M1 ;
        RECT 27.904 4.836 27.936 10.368 ;
  LAYER M2 ;
        RECT 22.444 10.252 27.956 10.284 ;
  LAYER M2 ;
        RECT 22.444 10.188 27.956 10.22 ;
  LAYER M2 ;
        RECT 22.444 10.124 27.956 10.156 ;
  LAYER M2 ;
        RECT 22.444 10.06 27.956 10.092 ;
  LAYER M2 ;
        RECT 22.444 9.996 27.956 10.028 ;
  LAYER M2 ;
        RECT 22.444 9.932 27.956 9.964 ;
  LAYER M2 ;
        RECT 22.444 9.868 27.956 9.9 ;
  LAYER M2 ;
        RECT 22.444 9.804 27.956 9.836 ;
  LAYER M2 ;
        RECT 22.444 9.74 27.956 9.772 ;
  LAYER M2 ;
        RECT 22.444 9.676 27.956 9.708 ;
  LAYER M2 ;
        RECT 22.444 9.612 27.956 9.644 ;
  LAYER M2 ;
        RECT 22.444 9.548 27.956 9.58 ;
  LAYER M2 ;
        RECT 22.444 9.484 27.956 9.516 ;
  LAYER M2 ;
        RECT 22.444 9.42 27.956 9.452 ;
  LAYER M2 ;
        RECT 22.444 9.356 27.956 9.388 ;
  LAYER M2 ;
        RECT 22.444 9.292 27.956 9.324 ;
  LAYER M2 ;
        RECT 22.444 9.228 27.956 9.26 ;
  LAYER M2 ;
        RECT 22.444 9.164 27.956 9.196 ;
  LAYER M2 ;
        RECT 22.444 9.1 27.956 9.132 ;
  LAYER M2 ;
        RECT 22.444 9.036 27.956 9.068 ;
  LAYER M2 ;
        RECT 22.444 8.972 27.956 9.004 ;
  LAYER M2 ;
        RECT 22.444 8.908 27.956 8.94 ;
  LAYER M2 ;
        RECT 22.444 8.844 27.956 8.876 ;
  LAYER M2 ;
        RECT 22.444 8.78 27.956 8.812 ;
  LAYER M2 ;
        RECT 22.444 8.716 27.956 8.748 ;
  LAYER M2 ;
        RECT 22.444 8.652 27.956 8.684 ;
  LAYER M2 ;
        RECT 22.444 8.588 27.956 8.62 ;
  LAYER M2 ;
        RECT 22.444 8.524 27.956 8.556 ;
  LAYER M2 ;
        RECT 22.444 8.46 27.956 8.492 ;
  LAYER M2 ;
        RECT 22.444 8.396 27.956 8.428 ;
  LAYER M2 ;
        RECT 22.444 8.332 27.956 8.364 ;
  LAYER M2 ;
        RECT 22.444 8.268 27.956 8.3 ;
  LAYER M2 ;
        RECT 22.444 8.204 27.956 8.236 ;
  LAYER M2 ;
        RECT 22.444 8.14 27.956 8.172 ;
  LAYER M2 ;
        RECT 22.444 8.076 27.956 8.108 ;
  LAYER M2 ;
        RECT 22.444 8.012 27.956 8.044 ;
  LAYER M2 ;
        RECT 22.444 7.948 27.956 7.98 ;
  LAYER M2 ;
        RECT 22.444 7.884 27.956 7.916 ;
  LAYER M2 ;
        RECT 22.444 7.82 27.956 7.852 ;
  LAYER M2 ;
        RECT 22.444 7.756 27.956 7.788 ;
  LAYER M2 ;
        RECT 22.444 7.692 27.956 7.724 ;
  LAYER M2 ;
        RECT 22.444 7.628 27.956 7.66 ;
  LAYER M2 ;
        RECT 22.444 7.564 27.956 7.596 ;
  LAYER M2 ;
        RECT 22.444 7.5 27.956 7.532 ;
  LAYER M2 ;
        RECT 22.444 7.436 27.956 7.468 ;
  LAYER M2 ;
        RECT 22.444 7.372 27.956 7.404 ;
  LAYER M2 ;
        RECT 22.444 7.308 27.956 7.34 ;
  LAYER M2 ;
        RECT 22.444 7.244 27.956 7.276 ;
  LAYER M2 ;
        RECT 22.444 7.18 27.956 7.212 ;
  LAYER M2 ;
        RECT 22.444 7.116 27.956 7.148 ;
  LAYER M2 ;
        RECT 22.444 7.052 27.956 7.084 ;
  LAYER M2 ;
        RECT 22.444 6.988 27.956 7.02 ;
  LAYER M2 ;
        RECT 22.444 6.924 27.956 6.956 ;
  LAYER M2 ;
        RECT 22.444 6.86 27.956 6.892 ;
  LAYER M2 ;
        RECT 22.444 6.796 27.956 6.828 ;
  LAYER M2 ;
        RECT 22.444 6.732 27.956 6.764 ;
  LAYER M2 ;
        RECT 22.444 6.668 27.956 6.7 ;
  LAYER M2 ;
        RECT 22.444 6.604 27.956 6.636 ;
  LAYER M2 ;
        RECT 22.444 6.54 27.956 6.572 ;
  LAYER M2 ;
        RECT 22.444 6.476 27.956 6.508 ;
  LAYER M2 ;
        RECT 22.444 6.412 27.956 6.444 ;
  LAYER M2 ;
        RECT 22.444 6.348 27.956 6.38 ;
  LAYER M2 ;
        RECT 22.444 6.284 27.956 6.316 ;
  LAYER M2 ;
        RECT 22.444 6.22 27.956 6.252 ;
  LAYER M2 ;
        RECT 22.444 6.156 27.956 6.188 ;
  LAYER M2 ;
        RECT 22.444 6.092 27.956 6.124 ;
  LAYER M2 ;
        RECT 22.444 6.028 27.956 6.06 ;
  LAYER M2 ;
        RECT 22.444 5.964 27.956 5.996 ;
  LAYER M2 ;
        RECT 22.444 5.9 27.956 5.932 ;
  LAYER M2 ;
        RECT 22.444 5.836 27.956 5.868 ;
  LAYER M2 ;
        RECT 22.444 5.772 27.956 5.804 ;
  LAYER M2 ;
        RECT 22.444 5.708 27.956 5.74 ;
  LAYER M2 ;
        RECT 22.444 5.644 27.956 5.676 ;
  LAYER M2 ;
        RECT 22.444 5.58 27.956 5.612 ;
  LAYER M2 ;
        RECT 22.444 5.516 27.956 5.548 ;
  LAYER M2 ;
        RECT 22.444 5.452 27.956 5.484 ;
  LAYER M2 ;
        RECT 22.444 5.388 27.956 5.42 ;
  LAYER M2 ;
        RECT 22.444 5.324 27.956 5.356 ;
  LAYER M2 ;
        RECT 22.444 5.26 27.956 5.292 ;
  LAYER M2 ;
        RECT 22.444 5.196 27.956 5.228 ;
  LAYER M2 ;
        RECT 22.444 5.132 27.956 5.164 ;
  LAYER M2 ;
        RECT 22.444 5.068 27.956 5.1 ;
  LAYER M2 ;
        RECT 22.444 5.004 27.956 5.036 ;
  LAYER M2 ;
        RECT 22.444 4.94 27.956 4.972 ;
  LAYER M3 ;
        RECT 22.464 4.836 22.496 10.368 ;
  LAYER M3 ;
        RECT 22.528 4.836 22.56 10.368 ;
  LAYER M3 ;
        RECT 22.592 4.836 22.624 10.368 ;
  LAYER M3 ;
        RECT 22.656 4.836 22.688 10.368 ;
  LAYER M3 ;
        RECT 22.72 4.836 22.752 10.368 ;
  LAYER M3 ;
        RECT 22.784 4.836 22.816 10.368 ;
  LAYER M3 ;
        RECT 22.848 4.836 22.88 10.368 ;
  LAYER M3 ;
        RECT 22.912 4.836 22.944 10.368 ;
  LAYER M3 ;
        RECT 22.976 4.836 23.008 10.368 ;
  LAYER M3 ;
        RECT 23.04 4.836 23.072 10.368 ;
  LAYER M3 ;
        RECT 23.104 4.836 23.136 10.368 ;
  LAYER M3 ;
        RECT 23.168 4.836 23.2 10.368 ;
  LAYER M3 ;
        RECT 23.232 4.836 23.264 10.368 ;
  LAYER M3 ;
        RECT 23.296 4.836 23.328 10.368 ;
  LAYER M3 ;
        RECT 23.36 4.836 23.392 10.368 ;
  LAYER M3 ;
        RECT 23.424 4.836 23.456 10.368 ;
  LAYER M3 ;
        RECT 23.488 4.836 23.52 10.368 ;
  LAYER M3 ;
        RECT 23.552 4.836 23.584 10.368 ;
  LAYER M3 ;
        RECT 23.616 4.836 23.648 10.368 ;
  LAYER M3 ;
        RECT 23.68 4.836 23.712 10.368 ;
  LAYER M3 ;
        RECT 23.744 4.836 23.776 10.368 ;
  LAYER M3 ;
        RECT 23.808 4.836 23.84 10.368 ;
  LAYER M3 ;
        RECT 23.872 4.836 23.904 10.368 ;
  LAYER M3 ;
        RECT 23.936 4.836 23.968 10.368 ;
  LAYER M3 ;
        RECT 24 4.836 24.032 10.368 ;
  LAYER M3 ;
        RECT 24.064 4.836 24.096 10.368 ;
  LAYER M3 ;
        RECT 24.128 4.836 24.16 10.368 ;
  LAYER M3 ;
        RECT 24.192 4.836 24.224 10.368 ;
  LAYER M3 ;
        RECT 24.256 4.836 24.288 10.368 ;
  LAYER M3 ;
        RECT 24.32 4.836 24.352 10.368 ;
  LAYER M3 ;
        RECT 24.384 4.836 24.416 10.368 ;
  LAYER M3 ;
        RECT 24.448 4.836 24.48 10.368 ;
  LAYER M3 ;
        RECT 24.512 4.836 24.544 10.368 ;
  LAYER M3 ;
        RECT 24.576 4.836 24.608 10.368 ;
  LAYER M3 ;
        RECT 24.64 4.836 24.672 10.368 ;
  LAYER M3 ;
        RECT 24.704 4.836 24.736 10.368 ;
  LAYER M3 ;
        RECT 24.768 4.836 24.8 10.368 ;
  LAYER M3 ;
        RECT 24.832 4.836 24.864 10.368 ;
  LAYER M3 ;
        RECT 24.896 4.836 24.928 10.368 ;
  LAYER M3 ;
        RECT 24.96 4.836 24.992 10.368 ;
  LAYER M3 ;
        RECT 25.024 4.836 25.056 10.368 ;
  LAYER M3 ;
        RECT 25.088 4.836 25.12 10.368 ;
  LAYER M3 ;
        RECT 25.152 4.836 25.184 10.368 ;
  LAYER M3 ;
        RECT 25.216 4.836 25.248 10.368 ;
  LAYER M3 ;
        RECT 25.28 4.836 25.312 10.368 ;
  LAYER M3 ;
        RECT 25.344 4.836 25.376 10.368 ;
  LAYER M3 ;
        RECT 25.408 4.836 25.44 10.368 ;
  LAYER M3 ;
        RECT 25.472 4.836 25.504 10.368 ;
  LAYER M3 ;
        RECT 25.536 4.836 25.568 10.368 ;
  LAYER M3 ;
        RECT 25.6 4.836 25.632 10.368 ;
  LAYER M3 ;
        RECT 25.664 4.836 25.696 10.368 ;
  LAYER M3 ;
        RECT 25.728 4.836 25.76 10.368 ;
  LAYER M3 ;
        RECT 25.792 4.836 25.824 10.368 ;
  LAYER M3 ;
        RECT 25.856 4.836 25.888 10.368 ;
  LAYER M3 ;
        RECT 25.92 4.836 25.952 10.368 ;
  LAYER M3 ;
        RECT 25.984 4.836 26.016 10.368 ;
  LAYER M3 ;
        RECT 26.048 4.836 26.08 10.368 ;
  LAYER M3 ;
        RECT 26.112 4.836 26.144 10.368 ;
  LAYER M3 ;
        RECT 26.176 4.836 26.208 10.368 ;
  LAYER M3 ;
        RECT 26.24 4.836 26.272 10.368 ;
  LAYER M3 ;
        RECT 26.304 4.836 26.336 10.368 ;
  LAYER M3 ;
        RECT 26.368 4.836 26.4 10.368 ;
  LAYER M3 ;
        RECT 26.432 4.836 26.464 10.368 ;
  LAYER M3 ;
        RECT 26.496 4.836 26.528 10.368 ;
  LAYER M3 ;
        RECT 26.56 4.836 26.592 10.368 ;
  LAYER M3 ;
        RECT 26.624 4.836 26.656 10.368 ;
  LAYER M3 ;
        RECT 26.688 4.836 26.72 10.368 ;
  LAYER M3 ;
        RECT 26.752 4.836 26.784 10.368 ;
  LAYER M3 ;
        RECT 26.816 4.836 26.848 10.368 ;
  LAYER M3 ;
        RECT 26.88 4.836 26.912 10.368 ;
  LAYER M3 ;
        RECT 26.944 4.836 26.976 10.368 ;
  LAYER M3 ;
        RECT 27.008 4.836 27.04 10.368 ;
  LAYER M3 ;
        RECT 27.072 4.836 27.104 10.368 ;
  LAYER M3 ;
        RECT 27.136 4.836 27.168 10.368 ;
  LAYER M3 ;
        RECT 27.2 4.836 27.232 10.368 ;
  LAYER M3 ;
        RECT 27.264 4.836 27.296 10.368 ;
  LAYER M3 ;
        RECT 27.328 4.836 27.36 10.368 ;
  LAYER M3 ;
        RECT 27.392 4.836 27.424 10.368 ;
  LAYER M3 ;
        RECT 27.456 4.836 27.488 10.368 ;
  LAYER M3 ;
        RECT 27.52 4.836 27.552 10.368 ;
  LAYER M3 ;
        RECT 27.584 4.836 27.616 10.368 ;
  LAYER M3 ;
        RECT 27.648 4.836 27.68 10.368 ;
  LAYER M3 ;
        RECT 27.712 4.836 27.744 10.368 ;
  LAYER M3 ;
        RECT 27.776 4.836 27.808 10.368 ;
  LAYER M3 ;
        RECT 27.84 4.836 27.872 10.368 ;
  LAYER M3 ;
        RECT 27.9 4.836 27.94 10.368 ;
  LAYER M2 ;
        RECT 22.204 4.856 28.196 4.888 ;
  LAYER M2 ;
        RECT 22.204 10.316 28.196 10.348 ;
  LAYER M1 ;
        RECT 28.224 12.9 28.256 13.644 ;
  LAYER M1 ;
        RECT 28.224 13.74 28.256 13.98 ;
  LAYER M1 ;
        RECT 28.224 14.496 28.256 14.736 ;
  LAYER M1 ;
        RECT 28.304 12.9 28.336 13.644 ;
  LAYER M1 ;
        RECT 28.144 12.9 28.176 13.644 ;
  LAYER M2 ;
        RECT 28.204 14.6 28.436 14.632 ;
  LAYER M2 ;
        RECT 28.204 12.92 28.436 12.952 ;
  LAYER M2 ;
        RECT 28.204 13.76 28.436 13.792 ;
  LAYER M2 ;
        RECT 28.124 13.004 28.356 13.036 ;
  LAYER M1 ;
        RECT 30.304 12.9 30.336 13.644 ;
  LAYER M1 ;
        RECT 30.304 13.74 30.336 13.98 ;
  LAYER M1 ;
        RECT 30.304 14.496 30.336 14.736 ;
  LAYER M1 ;
        RECT 30.224 12.9 30.256 13.644 ;
  LAYER M1 ;
        RECT 30.384 12.9 30.416 13.644 ;
  LAYER M2 ;
        RECT 30.124 14.6 30.356 14.632 ;
  LAYER M2 ;
        RECT 30.124 12.92 30.356 12.952 ;
  LAYER M2 ;
        RECT 30.124 13.76 30.356 13.792 ;
  LAYER M2 ;
        RECT 30.204 13.004 30.436 13.036 ;
  LAYER M1 ;
        RECT 29.984 6.264 30.016 7.008 ;
  LAYER M1 ;
        RECT 29.984 5.928 30.016 6.168 ;
  LAYER M1 ;
        RECT 29.984 5.172 30.016 5.412 ;
  LAYER M1 ;
        RECT 29.904 6.264 29.936 7.008 ;
  LAYER M1 ;
        RECT 30.064 6.264 30.096 7.008 ;
  LAYER M2 ;
        RECT 29.804 5.276 30.036 5.308 ;
  LAYER M2 ;
        RECT 29.804 6.956 30.036 6.988 ;
  LAYER M2 ;
        RECT 29.804 6.116 30.036 6.148 ;
  LAYER M2 ;
        RECT 29.884 6.872 30.116 6.904 ;
  LAYER M1 ;
        RECT 28.544 6.264 28.576 7.008 ;
  LAYER M1 ;
        RECT 28.544 5.928 28.576 6.168 ;
  LAYER M1 ;
        RECT 28.544 5.172 28.576 5.412 ;
  LAYER M1 ;
        RECT 28.624 6.264 28.656 7.008 ;
  LAYER M1 ;
        RECT 28.464 6.264 28.496 7.008 ;
  LAYER M2 ;
        RECT 28.524 5.276 28.756 5.308 ;
  LAYER M2 ;
        RECT 28.524 6.956 28.756 6.988 ;
  LAYER M2 ;
        RECT 28.524 6.116 28.756 6.148 ;
  LAYER M2 ;
        RECT 28.444 6.872 28.676 6.904 ;
  END 
END SWITCHED_CAPACITOR_FILTER
