MACRO CMC_S_NMOS_B_94218540_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CMC_S_NMOS_B_94218540_X1_Y1 0 0 ;
  SIZE 1280 BY 2352 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 1748 996 1780 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 68 516 100 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 764 152 996 184 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284 908 996 940 ;
    END
  END G
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204 236 436 268 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 844 320 1076 352 ;
    END
  END SB
  OBS
    LAYER M1 ;
      RECT 304 48 336 792 ;
    LAYER M1 ;
      RECT 304 888 336 1128 ;
    LAYER M1 ;
      RECT 304 1644 336 1884 ;
    LAYER M1 ;
      RECT 224 48 256 792 ;
    LAYER M1 ;
      RECT 384 48 416 792 ;
    LAYER M1 ;
      RECT 944 48 976 792 ;
    LAYER M1 ;
      RECT 944 888 976 1128 ;
    LAYER M1 ;
      RECT 944 1644 976 1884 ;
    LAYER M1 ;
      RECT 864 48 896 792 ;
    LAYER M1 ;
      RECT 1024 48 1056 792 ;
    LAYER V1 ;
      RECT 304 68 336 100 ;
    LAYER V1 ;
      RECT 304 908 336 940 ;
    LAYER V1 ;
      RECT 304 1748 336 1780 ;
    LAYER V1 ;
      RECT 944 152 976 184 ;
    LAYER V1 ;
      RECT 944 908 976 940 ;
    LAYER V1 ;
      RECT 944 1748 976 1780 ;
    LAYER V1 ;
      RECT 224 236 256 268 ;
    LAYER V1 ;
      RECT 384 236 416 268 ;
    LAYER V1 ;
      RECT 864 320 896 352 ;
    LAYER V1 ;
      RECT 1024 320 1056 352 ;
    LAYER V0 ;
      RECT 304 461 336 493 ;
    LAYER V0 ;
      RECT 304 545 336 577 ;
    LAYER V0 ;
      RECT 304 908 336 940 ;
    LAYER V0 ;
      RECT 304 1748 336 1780 ;
    LAYER V0 ;
      RECT 224 461 256 493 ;
    LAYER V0 ;
      RECT 224 545 256 577 ;
    LAYER V0 ;
      RECT 384 461 416 493 ;
    LAYER V0 ;
      RECT 384 545 416 577 ;
    LAYER V0 ;
      RECT 944 461 976 493 ;
    LAYER V0 ;
      RECT 944 545 976 577 ;
    LAYER V0 ;
      RECT 944 908 976 940 ;
    LAYER V0 ;
      RECT 944 1748 976 1780 ;
    LAYER V0 ;
      RECT 864 461 896 493 ;
    LAYER V0 ;
      RECT 864 545 896 577 ;
    LAYER V0 ;
      RECT 1024 461 1056 493 ;
    LAYER V0 ;
      RECT 1024 545 1056 577 ;
  END
END CMC_S_NMOS_B_94218540_X1_Y1
